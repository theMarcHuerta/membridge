/* Machine-generated using Migen */
module AccessArbitration(

);



endmodule
