/* Machine-generated using Migen */
module top(
	input clk,
	input rst,
	input [31:0] addr,
	input [63:0] data_in,
	input mem_write,
	input mem_read,
	output reg [63:0] data_out,
	output reg ready,
	input sys_clk,
	input sys_rst
);

reg [3:0] mem_ctrl_cmd_decoded = 4'd0;
reg [31:0] mem_ctrl_address = 32'd0;
reg [31:0] mem_ctrl_timer = 32'd0;
reg [1:0] mem_ctrl_state = 2'd0;
reg [63:0] mem_ctrl_memorycontroller0 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller2 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller3 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller4 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller5 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller6 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller7 = 64'd0;
reg [2:0] mem_ctrl_buffer_index = 3'd0;
reg [1:0] mem_ctrl_power_state = 2'd0;
reg [63:0] mem_ctrl_memorycontroller8 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller9 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller10 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller11 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller12 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller13 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller14 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller15 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller16 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller17 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller18 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller19 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller20 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller21 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller22 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller23 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller24 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller25 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller26 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller27 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller28 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller29 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller30 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller31 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller32 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller33 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller34 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller35 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller36 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller37 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller38 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller39 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller40 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller41 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller42 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller43 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller44 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller45 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller46 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller47 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller48 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller49 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller50 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller51 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller52 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller53 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller54 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller55 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller56 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller57 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller58 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller59 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller60 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller61 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller62 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller63 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller64 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller65 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller66 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller67 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller68 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller69 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller70 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller71 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller72 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller73 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller74 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller75 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller76 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller77 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller78 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller79 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller80 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller81 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller82 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller83 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller84 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller85 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller86 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller87 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller88 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller89 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller90 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller91 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller92 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller93 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller94 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller95 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller96 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller97 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller98 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller99 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller100 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller101 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller102 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller103 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller104 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller105 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller106 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller107 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller108 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller109 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller110 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller111 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller112 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller113 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller114 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller115 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller116 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller117 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller118 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller119 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller120 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller121 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller122 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller123 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller124 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller125 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller126 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller127 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller128 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller129 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller130 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller131 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller132 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller133 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller134 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller135 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller136 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller137 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller138 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller139 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller140 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller141 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller142 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller143 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller144 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller145 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller146 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller147 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller148 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller149 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller150 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller151 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller152 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller153 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller154 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller155 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller156 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller157 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller158 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller159 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller160 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller161 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller162 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller163 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller164 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller165 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller166 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller167 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller168 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller169 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller170 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller171 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller172 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller173 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller174 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller175 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller176 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller177 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller178 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller179 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller180 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller181 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller182 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller183 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller184 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller185 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller186 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller187 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller188 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller189 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller190 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller191 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller192 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller193 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller194 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller195 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller196 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller197 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller198 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller199 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller200 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller201 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller202 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller203 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller204 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller205 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller206 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller207 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller208 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller209 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller210 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller211 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller212 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller213 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller214 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller215 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller216 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller217 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller218 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller219 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller220 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller221 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller222 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller223 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller224 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller225 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller226 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller227 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller228 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller229 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller230 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller231 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller232 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller233 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller234 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller235 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller236 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller237 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller238 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller239 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller240 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller241 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller242 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller243 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller244 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller245 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller246 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller247 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller248 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller249 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller250 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller251 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller252 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller253 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller254 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller255 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller256 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller257 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller258 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller259 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller260 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller261 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller262 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller263 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller264 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller265 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller266 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller267 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller268 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller269 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller270 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller271 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller272 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller273 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller274 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller275 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller276 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller277 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller278 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller279 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller280 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller281 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller282 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller283 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller284 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller285 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller286 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller287 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller288 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller289 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller290 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller291 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller292 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller293 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller294 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller295 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller296 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller297 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller298 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller299 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller300 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller301 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller302 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller303 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller304 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller305 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller306 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller307 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller308 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller309 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller310 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller311 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller312 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller313 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller314 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller315 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller316 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller317 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller318 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller319 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller320 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller321 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller322 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller323 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller324 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller325 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller326 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller327 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller328 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller329 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller330 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller331 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller332 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller333 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller334 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller335 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller336 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller337 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller338 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller339 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller340 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller341 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller342 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller343 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller344 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller345 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller346 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller347 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller348 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller349 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller350 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller351 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller352 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller353 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller354 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller355 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller356 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller357 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller358 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller359 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller360 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller361 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller362 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller363 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller364 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller365 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller366 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller367 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller368 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller369 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller370 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller371 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller372 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller373 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller374 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller375 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller376 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller377 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller378 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller379 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller380 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller381 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller382 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller383 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller384 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller385 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller386 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller387 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller388 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller389 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller390 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller391 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller392 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller393 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller394 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller395 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller396 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller397 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller398 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller399 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller400 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller401 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller402 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller403 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller404 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller405 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller406 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller407 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller408 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller409 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller410 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller411 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller412 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller413 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller414 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller415 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller416 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller417 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller418 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller419 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller420 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller421 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller422 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller423 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller424 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller425 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller426 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller427 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller428 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller429 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller430 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller431 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller432 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller433 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller434 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller435 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller436 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller437 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller438 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller439 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller440 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller441 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller442 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller443 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller444 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller445 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller446 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller447 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller448 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller449 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller450 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller451 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller452 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller453 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller454 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller455 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller456 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller457 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller458 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller459 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller460 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller461 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller462 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller463 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller464 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller465 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller466 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller467 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller468 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller469 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller470 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller471 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller472 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller473 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller474 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller475 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller476 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller477 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller478 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller479 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller480 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller481 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller482 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller483 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller484 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller485 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller486 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller487 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller488 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller489 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller490 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller491 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller492 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller493 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller494 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller495 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller496 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller497 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller498 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller499 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller500 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller501 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller502 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller503 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller504 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller505 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller506 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller507 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller508 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller509 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller510 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller511 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller512 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller513 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller514 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller515 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller516 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller517 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller518 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller519 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller520 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller521 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller522 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller523 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller524 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller525 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller526 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller527 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller528 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller529 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller530 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller531 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller532 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller533 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller534 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller535 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller536 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller537 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller538 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller539 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller540 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller541 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller542 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller543 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller544 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller545 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller546 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller547 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller548 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller549 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller550 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller551 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller552 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller553 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller554 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller555 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller556 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller557 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller558 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller559 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller560 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller561 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller562 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller563 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller564 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller565 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller566 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller567 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller568 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller569 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller570 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller571 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller572 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller573 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller574 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller575 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller576 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller577 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller578 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller579 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller580 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller581 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller582 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller583 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller584 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller585 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller586 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller587 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller588 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller589 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller590 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller591 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller592 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller593 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller594 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller595 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller596 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller597 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller598 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller599 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller600 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller601 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller602 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller603 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller604 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller605 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller606 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller607 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller608 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller609 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller610 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller611 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller612 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller613 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller614 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller615 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller616 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller617 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller618 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller619 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller620 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller621 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller622 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller623 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller624 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller625 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller626 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller627 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller628 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller629 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller630 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller631 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller632 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller633 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller634 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller635 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller636 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller637 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller638 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller639 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller640 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller641 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller642 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller643 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller644 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller645 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller646 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller647 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller648 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller649 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller650 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller651 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller652 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller653 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller654 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller655 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller656 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller657 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller658 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller659 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller660 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller661 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller662 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller663 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller664 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller665 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller666 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller667 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller668 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller669 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller670 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller671 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller672 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller673 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller674 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller675 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller676 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller677 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller678 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller679 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller680 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller681 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller682 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller683 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller684 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller685 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller686 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller687 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller688 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller689 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller690 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller691 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller692 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller693 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller694 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller695 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller696 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller697 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller698 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller699 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller700 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller701 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller702 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller703 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller704 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller705 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller706 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller707 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller708 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller709 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller710 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller711 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller712 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller713 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller714 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller715 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller716 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller717 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller718 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller719 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller720 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller721 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller722 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller723 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller724 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller725 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller726 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller727 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller728 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller729 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller730 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller731 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller732 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller733 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller734 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller735 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller736 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller737 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller738 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller739 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller740 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller741 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller742 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller743 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller744 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller745 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller746 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller747 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller748 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller749 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller750 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller751 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller752 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller753 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller754 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller755 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller756 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller757 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller758 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller759 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller760 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller761 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller762 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller763 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller764 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller765 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller766 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller767 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller768 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller769 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller770 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller771 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller772 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller773 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller774 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller775 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller776 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller777 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller778 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller779 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller780 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller781 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller782 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller783 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller784 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller785 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller786 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller787 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller788 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller789 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller790 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller791 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller792 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller793 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller794 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller795 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller796 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller797 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller798 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller799 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller800 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller801 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller802 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller803 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller804 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller805 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller806 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller807 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller808 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller809 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller810 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller811 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller812 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller813 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller814 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller815 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller816 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller817 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller818 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller819 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller820 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller821 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller822 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller823 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller824 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller825 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller826 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller827 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller828 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller829 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller830 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller831 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller832 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller833 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller834 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller835 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller836 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller837 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller838 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller839 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller840 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller841 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller842 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller843 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller844 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller845 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller846 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller847 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller848 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller849 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller850 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller851 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller852 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller853 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller854 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller855 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller856 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller857 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller858 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller859 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller860 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller861 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller862 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller863 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller864 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller865 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller866 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller867 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller868 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller869 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller870 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller871 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller872 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller873 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller874 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller875 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller876 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller877 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller878 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller879 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller880 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller881 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller882 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller883 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller884 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller885 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller886 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller887 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller888 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller889 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller890 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller891 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller892 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller893 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller894 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller895 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller896 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller897 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller898 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller899 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller900 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller901 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller902 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller903 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller904 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller905 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller906 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller907 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller908 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller909 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller910 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller911 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller912 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller913 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller914 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller915 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller916 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller917 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller918 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller919 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller920 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller921 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller922 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller923 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller924 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller925 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller926 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller927 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller928 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller929 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller930 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller931 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller932 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller933 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller934 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller935 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller936 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller937 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller938 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller939 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller940 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller941 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller942 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller943 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller944 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller945 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller946 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller947 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller948 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller949 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller950 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller951 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller952 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller953 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller954 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller955 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller956 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller957 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller958 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller959 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller960 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller961 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller962 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller963 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller964 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller965 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller966 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller967 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller968 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller969 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller970 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller971 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller972 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller973 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller974 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller975 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller976 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller977 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller978 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller979 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller980 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller981 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller982 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller983 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller984 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller985 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller986 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller987 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller988 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller989 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller990 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller991 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller992 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller993 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller994 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller995 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller996 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller997 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller998 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller999 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1000 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1001 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1002 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1003 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1004 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1005 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1006 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1007 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1008 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1009 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1010 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1011 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1012 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1013 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1014 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1015 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1016 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1017 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1018 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1019 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1020 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1021 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1022 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1023 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1024 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1025 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1026 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1027 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1028 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1029 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1030 = 64'd0;
reg [63:0] mem_ctrl_memorycontroller1031 = 64'd0;
reg [63:0] verilog_output_t_lhs_array_muxed0 = 64'd0;
reg [63:0] verilog_output_f_rhs_array_muxed0;
reg [63:0] verilog_output_t_lhs_array_muxed1 = 64'd0;
reg [63:0] verilog_output_t_rhs_array_muxed;
reg [63:0] verilog_output_f_lhs_array_muxed = 64'd0;
reg [63:0] verilog_output_f_rhs_array_muxed1;

// synthesis translate_off
reg dummy_s;
initial dummy_s <= 1'd0;
// synthesis translate_on


// synthesis translate_off
reg dummy_d;
// synthesis translate_on
always @(*) begin
	verilog_output_f_rhs_array_muxed0 <= 64'd0;
	case (mem_ctrl_buffer_index)
		1'd0: begin
			verilog_output_f_rhs_array_muxed0 <= mem_ctrl_memorycontroller0;
		end
		1'd1: begin
			verilog_output_f_rhs_array_muxed0 <= mem_ctrl_memorycontroller1;
		end
		2'd2: begin
			verilog_output_f_rhs_array_muxed0 <= mem_ctrl_memorycontroller2;
		end
		2'd3: begin
			verilog_output_f_rhs_array_muxed0 <= mem_ctrl_memorycontroller3;
		end
		3'd4: begin
			verilog_output_f_rhs_array_muxed0 <= mem_ctrl_memorycontroller4;
		end
		3'd5: begin
			verilog_output_f_rhs_array_muxed0 <= mem_ctrl_memorycontroller5;
		end
		3'd6: begin
			verilog_output_f_rhs_array_muxed0 <= mem_ctrl_memorycontroller6;
		end
		default: begin
			verilog_output_f_rhs_array_muxed0 <= mem_ctrl_memorycontroller7;
		end
	endcase
// synthesis translate_off
	dummy_d <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_1;
// synthesis translate_on
always @(*) begin
	verilog_output_t_rhs_array_muxed <= 64'd0;
	case (mem_ctrl_address)
		1'd0: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller8;
		end
		1'd1: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller9;
		end
		2'd2: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller10;
		end
		2'd3: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller11;
		end
		3'd4: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller12;
		end
		3'd5: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller13;
		end
		3'd6: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller14;
		end
		3'd7: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller15;
		end
		4'd8: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller16;
		end
		4'd9: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller17;
		end
		4'd10: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller18;
		end
		4'd11: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller19;
		end
		4'd12: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller20;
		end
		4'd13: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller21;
		end
		4'd14: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller22;
		end
		4'd15: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller23;
		end
		5'd16: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller24;
		end
		5'd17: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller25;
		end
		5'd18: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller26;
		end
		5'd19: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller27;
		end
		5'd20: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller28;
		end
		5'd21: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller29;
		end
		5'd22: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller30;
		end
		5'd23: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller31;
		end
		5'd24: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller32;
		end
		5'd25: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller33;
		end
		5'd26: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller34;
		end
		5'd27: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller35;
		end
		5'd28: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller36;
		end
		5'd29: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller37;
		end
		5'd30: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller38;
		end
		5'd31: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller39;
		end
		6'd32: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller40;
		end
		6'd33: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller41;
		end
		6'd34: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller42;
		end
		6'd35: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller43;
		end
		6'd36: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller44;
		end
		6'd37: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller45;
		end
		6'd38: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller46;
		end
		6'd39: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller47;
		end
		6'd40: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller48;
		end
		6'd41: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller49;
		end
		6'd42: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller50;
		end
		6'd43: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller51;
		end
		6'd44: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller52;
		end
		6'd45: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller53;
		end
		6'd46: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller54;
		end
		6'd47: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller55;
		end
		6'd48: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller56;
		end
		6'd49: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller57;
		end
		6'd50: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller58;
		end
		6'd51: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller59;
		end
		6'd52: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller60;
		end
		6'd53: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller61;
		end
		6'd54: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller62;
		end
		6'd55: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller63;
		end
		6'd56: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller64;
		end
		6'd57: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller65;
		end
		6'd58: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller66;
		end
		6'd59: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller67;
		end
		6'd60: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller68;
		end
		6'd61: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller69;
		end
		6'd62: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller70;
		end
		6'd63: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller71;
		end
		7'd64: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller72;
		end
		7'd65: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller73;
		end
		7'd66: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller74;
		end
		7'd67: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller75;
		end
		7'd68: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller76;
		end
		7'd69: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller77;
		end
		7'd70: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller78;
		end
		7'd71: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller79;
		end
		7'd72: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller80;
		end
		7'd73: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller81;
		end
		7'd74: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller82;
		end
		7'd75: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller83;
		end
		7'd76: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller84;
		end
		7'd77: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller85;
		end
		7'd78: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller86;
		end
		7'd79: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller87;
		end
		7'd80: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller88;
		end
		7'd81: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller89;
		end
		7'd82: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller90;
		end
		7'd83: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller91;
		end
		7'd84: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller92;
		end
		7'd85: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller93;
		end
		7'd86: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller94;
		end
		7'd87: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller95;
		end
		7'd88: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller96;
		end
		7'd89: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller97;
		end
		7'd90: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller98;
		end
		7'd91: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller99;
		end
		7'd92: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller100;
		end
		7'd93: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller101;
		end
		7'd94: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller102;
		end
		7'd95: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller103;
		end
		7'd96: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller104;
		end
		7'd97: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller105;
		end
		7'd98: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller106;
		end
		7'd99: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller107;
		end
		7'd100: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller108;
		end
		7'd101: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller109;
		end
		7'd102: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller110;
		end
		7'd103: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller111;
		end
		7'd104: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller112;
		end
		7'd105: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller113;
		end
		7'd106: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller114;
		end
		7'd107: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller115;
		end
		7'd108: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller116;
		end
		7'd109: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller117;
		end
		7'd110: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller118;
		end
		7'd111: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller119;
		end
		7'd112: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller120;
		end
		7'd113: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller121;
		end
		7'd114: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller122;
		end
		7'd115: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller123;
		end
		7'd116: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller124;
		end
		7'd117: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller125;
		end
		7'd118: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller126;
		end
		7'd119: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller127;
		end
		7'd120: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller128;
		end
		7'd121: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller129;
		end
		7'd122: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller130;
		end
		7'd123: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller131;
		end
		7'd124: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller132;
		end
		7'd125: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller133;
		end
		7'd126: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller134;
		end
		7'd127: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller135;
		end
		8'd128: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller136;
		end
		8'd129: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller137;
		end
		8'd130: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller138;
		end
		8'd131: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller139;
		end
		8'd132: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller140;
		end
		8'd133: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller141;
		end
		8'd134: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller142;
		end
		8'd135: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller143;
		end
		8'd136: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller144;
		end
		8'd137: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller145;
		end
		8'd138: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller146;
		end
		8'd139: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller147;
		end
		8'd140: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller148;
		end
		8'd141: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller149;
		end
		8'd142: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller150;
		end
		8'd143: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller151;
		end
		8'd144: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller152;
		end
		8'd145: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller153;
		end
		8'd146: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller154;
		end
		8'd147: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller155;
		end
		8'd148: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller156;
		end
		8'd149: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller157;
		end
		8'd150: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller158;
		end
		8'd151: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller159;
		end
		8'd152: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller160;
		end
		8'd153: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller161;
		end
		8'd154: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller162;
		end
		8'd155: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller163;
		end
		8'd156: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller164;
		end
		8'd157: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller165;
		end
		8'd158: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller166;
		end
		8'd159: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller167;
		end
		8'd160: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller168;
		end
		8'd161: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller169;
		end
		8'd162: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller170;
		end
		8'd163: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller171;
		end
		8'd164: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller172;
		end
		8'd165: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller173;
		end
		8'd166: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller174;
		end
		8'd167: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller175;
		end
		8'd168: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller176;
		end
		8'd169: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller177;
		end
		8'd170: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller178;
		end
		8'd171: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller179;
		end
		8'd172: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller180;
		end
		8'd173: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller181;
		end
		8'd174: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller182;
		end
		8'd175: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller183;
		end
		8'd176: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller184;
		end
		8'd177: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller185;
		end
		8'd178: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller186;
		end
		8'd179: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller187;
		end
		8'd180: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller188;
		end
		8'd181: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller189;
		end
		8'd182: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller190;
		end
		8'd183: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller191;
		end
		8'd184: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller192;
		end
		8'd185: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller193;
		end
		8'd186: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller194;
		end
		8'd187: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller195;
		end
		8'd188: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller196;
		end
		8'd189: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller197;
		end
		8'd190: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller198;
		end
		8'd191: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller199;
		end
		8'd192: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller200;
		end
		8'd193: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller201;
		end
		8'd194: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller202;
		end
		8'd195: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller203;
		end
		8'd196: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller204;
		end
		8'd197: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller205;
		end
		8'd198: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller206;
		end
		8'd199: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller207;
		end
		8'd200: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller208;
		end
		8'd201: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller209;
		end
		8'd202: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller210;
		end
		8'd203: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller211;
		end
		8'd204: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller212;
		end
		8'd205: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller213;
		end
		8'd206: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller214;
		end
		8'd207: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller215;
		end
		8'd208: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller216;
		end
		8'd209: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller217;
		end
		8'd210: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller218;
		end
		8'd211: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller219;
		end
		8'd212: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller220;
		end
		8'd213: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller221;
		end
		8'd214: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller222;
		end
		8'd215: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller223;
		end
		8'd216: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller224;
		end
		8'd217: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller225;
		end
		8'd218: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller226;
		end
		8'd219: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller227;
		end
		8'd220: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller228;
		end
		8'd221: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller229;
		end
		8'd222: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller230;
		end
		8'd223: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller231;
		end
		8'd224: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller232;
		end
		8'd225: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller233;
		end
		8'd226: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller234;
		end
		8'd227: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller235;
		end
		8'd228: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller236;
		end
		8'd229: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller237;
		end
		8'd230: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller238;
		end
		8'd231: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller239;
		end
		8'd232: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller240;
		end
		8'd233: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller241;
		end
		8'd234: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller242;
		end
		8'd235: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller243;
		end
		8'd236: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller244;
		end
		8'd237: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller245;
		end
		8'd238: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller246;
		end
		8'd239: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller247;
		end
		8'd240: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller248;
		end
		8'd241: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller249;
		end
		8'd242: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller250;
		end
		8'd243: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller251;
		end
		8'd244: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller252;
		end
		8'd245: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller253;
		end
		8'd246: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller254;
		end
		8'd247: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller255;
		end
		8'd248: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller256;
		end
		8'd249: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller257;
		end
		8'd250: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller258;
		end
		8'd251: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller259;
		end
		8'd252: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller260;
		end
		8'd253: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller261;
		end
		8'd254: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller262;
		end
		8'd255: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller263;
		end
		9'd256: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller264;
		end
		9'd257: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller265;
		end
		9'd258: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller266;
		end
		9'd259: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller267;
		end
		9'd260: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller268;
		end
		9'd261: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller269;
		end
		9'd262: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller270;
		end
		9'd263: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller271;
		end
		9'd264: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller272;
		end
		9'd265: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller273;
		end
		9'd266: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller274;
		end
		9'd267: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller275;
		end
		9'd268: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller276;
		end
		9'd269: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller277;
		end
		9'd270: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller278;
		end
		9'd271: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller279;
		end
		9'd272: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller280;
		end
		9'd273: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller281;
		end
		9'd274: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller282;
		end
		9'd275: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller283;
		end
		9'd276: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller284;
		end
		9'd277: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller285;
		end
		9'd278: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller286;
		end
		9'd279: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller287;
		end
		9'd280: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller288;
		end
		9'd281: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller289;
		end
		9'd282: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller290;
		end
		9'd283: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller291;
		end
		9'd284: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller292;
		end
		9'd285: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller293;
		end
		9'd286: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller294;
		end
		9'd287: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller295;
		end
		9'd288: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller296;
		end
		9'd289: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller297;
		end
		9'd290: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller298;
		end
		9'd291: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller299;
		end
		9'd292: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller300;
		end
		9'd293: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller301;
		end
		9'd294: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller302;
		end
		9'd295: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller303;
		end
		9'd296: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller304;
		end
		9'd297: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller305;
		end
		9'd298: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller306;
		end
		9'd299: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller307;
		end
		9'd300: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller308;
		end
		9'd301: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller309;
		end
		9'd302: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller310;
		end
		9'd303: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller311;
		end
		9'd304: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller312;
		end
		9'd305: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller313;
		end
		9'd306: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller314;
		end
		9'd307: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller315;
		end
		9'd308: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller316;
		end
		9'd309: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller317;
		end
		9'd310: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller318;
		end
		9'd311: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller319;
		end
		9'd312: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller320;
		end
		9'd313: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller321;
		end
		9'd314: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller322;
		end
		9'd315: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller323;
		end
		9'd316: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller324;
		end
		9'd317: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller325;
		end
		9'd318: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller326;
		end
		9'd319: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller327;
		end
		9'd320: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller328;
		end
		9'd321: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller329;
		end
		9'd322: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller330;
		end
		9'd323: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller331;
		end
		9'd324: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller332;
		end
		9'd325: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller333;
		end
		9'd326: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller334;
		end
		9'd327: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller335;
		end
		9'd328: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller336;
		end
		9'd329: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller337;
		end
		9'd330: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller338;
		end
		9'd331: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller339;
		end
		9'd332: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller340;
		end
		9'd333: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller341;
		end
		9'd334: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller342;
		end
		9'd335: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller343;
		end
		9'd336: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller344;
		end
		9'd337: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller345;
		end
		9'd338: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller346;
		end
		9'd339: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller347;
		end
		9'd340: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller348;
		end
		9'd341: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller349;
		end
		9'd342: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller350;
		end
		9'd343: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller351;
		end
		9'd344: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller352;
		end
		9'd345: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller353;
		end
		9'd346: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller354;
		end
		9'd347: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller355;
		end
		9'd348: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller356;
		end
		9'd349: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller357;
		end
		9'd350: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller358;
		end
		9'd351: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller359;
		end
		9'd352: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller360;
		end
		9'd353: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller361;
		end
		9'd354: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller362;
		end
		9'd355: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller363;
		end
		9'd356: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller364;
		end
		9'd357: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller365;
		end
		9'd358: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller366;
		end
		9'd359: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller367;
		end
		9'd360: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller368;
		end
		9'd361: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller369;
		end
		9'd362: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller370;
		end
		9'd363: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller371;
		end
		9'd364: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller372;
		end
		9'd365: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller373;
		end
		9'd366: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller374;
		end
		9'd367: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller375;
		end
		9'd368: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller376;
		end
		9'd369: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller377;
		end
		9'd370: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller378;
		end
		9'd371: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller379;
		end
		9'd372: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller380;
		end
		9'd373: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller381;
		end
		9'd374: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller382;
		end
		9'd375: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller383;
		end
		9'd376: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller384;
		end
		9'd377: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller385;
		end
		9'd378: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller386;
		end
		9'd379: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller387;
		end
		9'd380: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller388;
		end
		9'd381: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller389;
		end
		9'd382: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller390;
		end
		9'd383: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller391;
		end
		9'd384: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller392;
		end
		9'd385: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller393;
		end
		9'd386: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller394;
		end
		9'd387: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller395;
		end
		9'd388: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller396;
		end
		9'd389: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller397;
		end
		9'd390: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller398;
		end
		9'd391: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller399;
		end
		9'd392: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller400;
		end
		9'd393: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller401;
		end
		9'd394: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller402;
		end
		9'd395: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller403;
		end
		9'd396: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller404;
		end
		9'd397: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller405;
		end
		9'd398: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller406;
		end
		9'd399: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller407;
		end
		9'd400: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller408;
		end
		9'd401: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller409;
		end
		9'd402: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller410;
		end
		9'd403: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller411;
		end
		9'd404: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller412;
		end
		9'd405: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller413;
		end
		9'd406: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller414;
		end
		9'd407: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller415;
		end
		9'd408: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller416;
		end
		9'd409: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller417;
		end
		9'd410: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller418;
		end
		9'd411: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller419;
		end
		9'd412: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller420;
		end
		9'd413: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller421;
		end
		9'd414: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller422;
		end
		9'd415: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller423;
		end
		9'd416: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller424;
		end
		9'd417: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller425;
		end
		9'd418: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller426;
		end
		9'd419: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller427;
		end
		9'd420: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller428;
		end
		9'd421: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller429;
		end
		9'd422: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller430;
		end
		9'd423: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller431;
		end
		9'd424: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller432;
		end
		9'd425: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller433;
		end
		9'd426: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller434;
		end
		9'd427: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller435;
		end
		9'd428: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller436;
		end
		9'd429: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller437;
		end
		9'd430: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller438;
		end
		9'd431: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller439;
		end
		9'd432: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller440;
		end
		9'd433: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller441;
		end
		9'd434: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller442;
		end
		9'd435: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller443;
		end
		9'd436: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller444;
		end
		9'd437: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller445;
		end
		9'd438: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller446;
		end
		9'd439: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller447;
		end
		9'd440: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller448;
		end
		9'd441: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller449;
		end
		9'd442: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller450;
		end
		9'd443: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller451;
		end
		9'd444: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller452;
		end
		9'd445: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller453;
		end
		9'd446: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller454;
		end
		9'd447: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller455;
		end
		9'd448: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller456;
		end
		9'd449: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller457;
		end
		9'd450: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller458;
		end
		9'd451: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller459;
		end
		9'd452: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller460;
		end
		9'd453: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller461;
		end
		9'd454: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller462;
		end
		9'd455: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller463;
		end
		9'd456: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller464;
		end
		9'd457: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller465;
		end
		9'd458: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller466;
		end
		9'd459: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller467;
		end
		9'd460: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller468;
		end
		9'd461: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller469;
		end
		9'd462: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller470;
		end
		9'd463: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller471;
		end
		9'd464: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller472;
		end
		9'd465: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller473;
		end
		9'd466: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller474;
		end
		9'd467: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller475;
		end
		9'd468: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller476;
		end
		9'd469: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller477;
		end
		9'd470: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller478;
		end
		9'd471: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller479;
		end
		9'd472: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller480;
		end
		9'd473: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller481;
		end
		9'd474: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller482;
		end
		9'd475: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller483;
		end
		9'd476: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller484;
		end
		9'd477: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller485;
		end
		9'd478: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller486;
		end
		9'd479: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller487;
		end
		9'd480: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller488;
		end
		9'd481: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller489;
		end
		9'd482: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller490;
		end
		9'd483: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller491;
		end
		9'd484: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller492;
		end
		9'd485: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller493;
		end
		9'd486: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller494;
		end
		9'd487: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller495;
		end
		9'd488: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller496;
		end
		9'd489: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller497;
		end
		9'd490: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller498;
		end
		9'd491: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller499;
		end
		9'd492: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller500;
		end
		9'd493: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller501;
		end
		9'd494: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller502;
		end
		9'd495: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller503;
		end
		9'd496: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller504;
		end
		9'd497: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller505;
		end
		9'd498: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller506;
		end
		9'd499: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller507;
		end
		9'd500: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller508;
		end
		9'd501: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller509;
		end
		9'd502: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller510;
		end
		9'd503: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller511;
		end
		9'd504: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller512;
		end
		9'd505: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller513;
		end
		9'd506: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller514;
		end
		9'd507: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller515;
		end
		9'd508: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller516;
		end
		9'd509: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller517;
		end
		9'd510: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller518;
		end
		9'd511: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller519;
		end
		10'd512: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller520;
		end
		10'd513: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller521;
		end
		10'd514: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller522;
		end
		10'd515: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller523;
		end
		10'd516: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller524;
		end
		10'd517: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller525;
		end
		10'd518: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller526;
		end
		10'd519: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller527;
		end
		10'd520: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller528;
		end
		10'd521: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller529;
		end
		10'd522: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller530;
		end
		10'd523: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller531;
		end
		10'd524: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller532;
		end
		10'd525: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller533;
		end
		10'd526: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller534;
		end
		10'd527: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller535;
		end
		10'd528: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller536;
		end
		10'd529: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller537;
		end
		10'd530: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller538;
		end
		10'd531: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller539;
		end
		10'd532: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller540;
		end
		10'd533: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller541;
		end
		10'd534: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller542;
		end
		10'd535: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller543;
		end
		10'd536: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller544;
		end
		10'd537: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller545;
		end
		10'd538: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller546;
		end
		10'd539: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller547;
		end
		10'd540: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller548;
		end
		10'd541: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller549;
		end
		10'd542: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller550;
		end
		10'd543: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller551;
		end
		10'd544: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller552;
		end
		10'd545: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller553;
		end
		10'd546: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller554;
		end
		10'd547: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller555;
		end
		10'd548: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller556;
		end
		10'd549: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller557;
		end
		10'd550: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller558;
		end
		10'd551: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller559;
		end
		10'd552: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller560;
		end
		10'd553: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller561;
		end
		10'd554: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller562;
		end
		10'd555: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller563;
		end
		10'd556: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller564;
		end
		10'd557: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller565;
		end
		10'd558: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller566;
		end
		10'd559: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller567;
		end
		10'd560: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller568;
		end
		10'd561: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller569;
		end
		10'd562: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller570;
		end
		10'd563: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller571;
		end
		10'd564: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller572;
		end
		10'd565: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller573;
		end
		10'd566: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller574;
		end
		10'd567: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller575;
		end
		10'd568: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller576;
		end
		10'd569: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller577;
		end
		10'd570: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller578;
		end
		10'd571: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller579;
		end
		10'd572: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller580;
		end
		10'd573: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller581;
		end
		10'd574: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller582;
		end
		10'd575: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller583;
		end
		10'd576: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller584;
		end
		10'd577: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller585;
		end
		10'd578: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller586;
		end
		10'd579: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller587;
		end
		10'd580: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller588;
		end
		10'd581: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller589;
		end
		10'd582: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller590;
		end
		10'd583: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller591;
		end
		10'd584: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller592;
		end
		10'd585: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller593;
		end
		10'd586: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller594;
		end
		10'd587: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller595;
		end
		10'd588: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller596;
		end
		10'd589: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller597;
		end
		10'd590: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller598;
		end
		10'd591: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller599;
		end
		10'd592: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller600;
		end
		10'd593: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller601;
		end
		10'd594: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller602;
		end
		10'd595: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller603;
		end
		10'd596: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller604;
		end
		10'd597: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller605;
		end
		10'd598: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller606;
		end
		10'd599: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller607;
		end
		10'd600: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller608;
		end
		10'd601: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller609;
		end
		10'd602: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller610;
		end
		10'd603: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller611;
		end
		10'd604: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller612;
		end
		10'd605: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller613;
		end
		10'd606: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller614;
		end
		10'd607: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller615;
		end
		10'd608: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller616;
		end
		10'd609: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller617;
		end
		10'd610: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller618;
		end
		10'd611: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller619;
		end
		10'd612: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller620;
		end
		10'd613: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller621;
		end
		10'd614: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller622;
		end
		10'd615: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller623;
		end
		10'd616: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller624;
		end
		10'd617: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller625;
		end
		10'd618: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller626;
		end
		10'd619: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller627;
		end
		10'd620: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller628;
		end
		10'd621: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller629;
		end
		10'd622: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller630;
		end
		10'd623: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller631;
		end
		10'd624: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller632;
		end
		10'd625: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller633;
		end
		10'd626: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller634;
		end
		10'd627: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller635;
		end
		10'd628: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller636;
		end
		10'd629: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller637;
		end
		10'd630: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller638;
		end
		10'd631: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller639;
		end
		10'd632: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller640;
		end
		10'd633: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller641;
		end
		10'd634: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller642;
		end
		10'd635: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller643;
		end
		10'd636: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller644;
		end
		10'd637: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller645;
		end
		10'd638: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller646;
		end
		10'd639: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller647;
		end
		10'd640: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller648;
		end
		10'd641: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller649;
		end
		10'd642: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller650;
		end
		10'd643: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller651;
		end
		10'd644: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller652;
		end
		10'd645: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller653;
		end
		10'd646: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller654;
		end
		10'd647: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller655;
		end
		10'd648: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller656;
		end
		10'd649: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller657;
		end
		10'd650: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller658;
		end
		10'd651: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller659;
		end
		10'd652: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller660;
		end
		10'd653: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller661;
		end
		10'd654: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller662;
		end
		10'd655: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller663;
		end
		10'd656: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller664;
		end
		10'd657: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller665;
		end
		10'd658: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller666;
		end
		10'd659: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller667;
		end
		10'd660: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller668;
		end
		10'd661: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller669;
		end
		10'd662: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller670;
		end
		10'd663: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller671;
		end
		10'd664: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller672;
		end
		10'd665: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller673;
		end
		10'd666: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller674;
		end
		10'd667: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller675;
		end
		10'd668: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller676;
		end
		10'd669: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller677;
		end
		10'd670: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller678;
		end
		10'd671: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller679;
		end
		10'd672: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller680;
		end
		10'd673: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller681;
		end
		10'd674: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller682;
		end
		10'd675: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller683;
		end
		10'd676: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller684;
		end
		10'd677: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller685;
		end
		10'd678: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller686;
		end
		10'd679: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller687;
		end
		10'd680: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller688;
		end
		10'd681: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller689;
		end
		10'd682: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller690;
		end
		10'd683: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller691;
		end
		10'd684: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller692;
		end
		10'd685: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller693;
		end
		10'd686: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller694;
		end
		10'd687: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller695;
		end
		10'd688: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller696;
		end
		10'd689: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller697;
		end
		10'd690: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller698;
		end
		10'd691: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller699;
		end
		10'd692: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller700;
		end
		10'd693: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller701;
		end
		10'd694: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller702;
		end
		10'd695: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller703;
		end
		10'd696: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller704;
		end
		10'd697: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller705;
		end
		10'd698: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller706;
		end
		10'd699: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller707;
		end
		10'd700: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller708;
		end
		10'd701: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller709;
		end
		10'd702: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller710;
		end
		10'd703: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller711;
		end
		10'd704: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller712;
		end
		10'd705: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller713;
		end
		10'd706: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller714;
		end
		10'd707: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller715;
		end
		10'd708: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller716;
		end
		10'd709: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller717;
		end
		10'd710: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller718;
		end
		10'd711: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller719;
		end
		10'd712: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller720;
		end
		10'd713: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller721;
		end
		10'd714: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller722;
		end
		10'd715: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller723;
		end
		10'd716: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller724;
		end
		10'd717: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller725;
		end
		10'd718: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller726;
		end
		10'd719: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller727;
		end
		10'd720: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller728;
		end
		10'd721: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller729;
		end
		10'd722: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller730;
		end
		10'd723: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller731;
		end
		10'd724: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller732;
		end
		10'd725: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller733;
		end
		10'd726: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller734;
		end
		10'd727: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller735;
		end
		10'd728: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller736;
		end
		10'd729: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller737;
		end
		10'd730: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller738;
		end
		10'd731: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller739;
		end
		10'd732: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller740;
		end
		10'd733: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller741;
		end
		10'd734: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller742;
		end
		10'd735: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller743;
		end
		10'd736: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller744;
		end
		10'd737: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller745;
		end
		10'd738: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller746;
		end
		10'd739: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller747;
		end
		10'd740: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller748;
		end
		10'd741: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller749;
		end
		10'd742: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller750;
		end
		10'd743: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller751;
		end
		10'd744: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller752;
		end
		10'd745: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller753;
		end
		10'd746: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller754;
		end
		10'd747: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller755;
		end
		10'd748: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller756;
		end
		10'd749: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller757;
		end
		10'd750: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller758;
		end
		10'd751: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller759;
		end
		10'd752: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller760;
		end
		10'd753: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller761;
		end
		10'd754: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller762;
		end
		10'd755: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller763;
		end
		10'd756: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller764;
		end
		10'd757: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller765;
		end
		10'd758: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller766;
		end
		10'd759: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller767;
		end
		10'd760: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller768;
		end
		10'd761: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller769;
		end
		10'd762: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller770;
		end
		10'd763: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller771;
		end
		10'd764: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller772;
		end
		10'd765: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller773;
		end
		10'd766: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller774;
		end
		10'd767: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller775;
		end
		10'd768: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller776;
		end
		10'd769: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller777;
		end
		10'd770: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller778;
		end
		10'd771: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller779;
		end
		10'd772: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller780;
		end
		10'd773: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller781;
		end
		10'd774: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller782;
		end
		10'd775: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller783;
		end
		10'd776: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller784;
		end
		10'd777: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller785;
		end
		10'd778: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller786;
		end
		10'd779: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller787;
		end
		10'd780: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller788;
		end
		10'd781: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller789;
		end
		10'd782: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller790;
		end
		10'd783: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller791;
		end
		10'd784: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller792;
		end
		10'd785: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller793;
		end
		10'd786: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller794;
		end
		10'd787: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller795;
		end
		10'd788: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller796;
		end
		10'd789: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller797;
		end
		10'd790: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller798;
		end
		10'd791: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller799;
		end
		10'd792: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller800;
		end
		10'd793: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller801;
		end
		10'd794: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller802;
		end
		10'd795: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller803;
		end
		10'd796: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller804;
		end
		10'd797: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller805;
		end
		10'd798: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller806;
		end
		10'd799: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller807;
		end
		10'd800: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller808;
		end
		10'd801: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller809;
		end
		10'd802: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller810;
		end
		10'd803: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller811;
		end
		10'd804: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller812;
		end
		10'd805: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller813;
		end
		10'd806: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller814;
		end
		10'd807: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller815;
		end
		10'd808: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller816;
		end
		10'd809: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller817;
		end
		10'd810: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller818;
		end
		10'd811: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller819;
		end
		10'd812: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller820;
		end
		10'd813: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller821;
		end
		10'd814: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller822;
		end
		10'd815: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller823;
		end
		10'd816: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller824;
		end
		10'd817: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller825;
		end
		10'd818: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller826;
		end
		10'd819: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller827;
		end
		10'd820: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller828;
		end
		10'd821: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller829;
		end
		10'd822: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller830;
		end
		10'd823: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller831;
		end
		10'd824: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller832;
		end
		10'd825: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller833;
		end
		10'd826: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller834;
		end
		10'd827: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller835;
		end
		10'd828: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller836;
		end
		10'd829: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller837;
		end
		10'd830: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller838;
		end
		10'd831: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller839;
		end
		10'd832: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller840;
		end
		10'd833: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller841;
		end
		10'd834: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller842;
		end
		10'd835: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller843;
		end
		10'd836: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller844;
		end
		10'd837: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller845;
		end
		10'd838: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller846;
		end
		10'd839: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller847;
		end
		10'd840: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller848;
		end
		10'd841: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller849;
		end
		10'd842: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller850;
		end
		10'd843: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller851;
		end
		10'd844: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller852;
		end
		10'd845: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller853;
		end
		10'd846: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller854;
		end
		10'd847: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller855;
		end
		10'd848: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller856;
		end
		10'd849: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller857;
		end
		10'd850: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller858;
		end
		10'd851: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller859;
		end
		10'd852: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller860;
		end
		10'd853: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller861;
		end
		10'd854: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller862;
		end
		10'd855: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller863;
		end
		10'd856: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller864;
		end
		10'd857: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller865;
		end
		10'd858: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller866;
		end
		10'd859: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller867;
		end
		10'd860: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller868;
		end
		10'd861: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller869;
		end
		10'd862: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller870;
		end
		10'd863: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller871;
		end
		10'd864: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller872;
		end
		10'd865: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller873;
		end
		10'd866: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller874;
		end
		10'd867: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller875;
		end
		10'd868: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller876;
		end
		10'd869: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller877;
		end
		10'd870: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller878;
		end
		10'd871: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller879;
		end
		10'd872: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller880;
		end
		10'd873: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller881;
		end
		10'd874: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller882;
		end
		10'd875: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller883;
		end
		10'd876: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller884;
		end
		10'd877: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller885;
		end
		10'd878: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller886;
		end
		10'd879: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller887;
		end
		10'd880: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller888;
		end
		10'd881: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller889;
		end
		10'd882: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller890;
		end
		10'd883: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller891;
		end
		10'd884: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller892;
		end
		10'd885: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller893;
		end
		10'd886: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller894;
		end
		10'd887: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller895;
		end
		10'd888: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller896;
		end
		10'd889: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller897;
		end
		10'd890: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller898;
		end
		10'd891: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller899;
		end
		10'd892: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller900;
		end
		10'd893: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller901;
		end
		10'd894: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller902;
		end
		10'd895: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller903;
		end
		10'd896: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller904;
		end
		10'd897: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller905;
		end
		10'd898: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller906;
		end
		10'd899: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller907;
		end
		10'd900: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller908;
		end
		10'd901: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller909;
		end
		10'd902: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller910;
		end
		10'd903: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller911;
		end
		10'd904: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller912;
		end
		10'd905: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller913;
		end
		10'd906: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller914;
		end
		10'd907: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller915;
		end
		10'd908: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller916;
		end
		10'd909: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller917;
		end
		10'd910: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller918;
		end
		10'd911: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller919;
		end
		10'd912: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller920;
		end
		10'd913: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller921;
		end
		10'd914: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller922;
		end
		10'd915: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller923;
		end
		10'd916: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller924;
		end
		10'd917: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller925;
		end
		10'd918: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller926;
		end
		10'd919: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller927;
		end
		10'd920: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller928;
		end
		10'd921: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller929;
		end
		10'd922: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller930;
		end
		10'd923: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller931;
		end
		10'd924: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller932;
		end
		10'd925: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller933;
		end
		10'd926: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller934;
		end
		10'd927: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller935;
		end
		10'd928: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller936;
		end
		10'd929: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller937;
		end
		10'd930: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller938;
		end
		10'd931: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller939;
		end
		10'd932: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller940;
		end
		10'd933: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller941;
		end
		10'd934: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller942;
		end
		10'd935: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller943;
		end
		10'd936: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller944;
		end
		10'd937: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller945;
		end
		10'd938: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller946;
		end
		10'd939: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller947;
		end
		10'd940: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller948;
		end
		10'd941: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller949;
		end
		10'd942: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller950;
		end
		10'd943: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller951;
		end
		10'd944: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller952;
		end
		10'd945: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller953;
		end
		10'd946: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller954;
		end
		10'd947: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller955;
		end
		10'd948: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller956;
		end
		10'd949: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller957;
		end
		10'd950: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller958;
		end
		10'd951: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller959;
		end
		10'd952: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller960;
		end
		10'd953: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller961;
		end
		10'd954: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller962;
		end
		10'd955: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller963;
		end
		10'd956: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller964;
		end
		10'd957: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller965;
		end
		10'd958: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller966;
		end
		10'd959: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller967;
		end
		10'd960: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller968;
		end
		10'd961: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller969;
		end
		10'd962: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller970;
		end
		10'd963: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller971;
		end
		10'd964: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller972;
		end
		10'd965: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller973;
		end
		10'd966: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller974;
		end
		10'd967: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller975;
		end
		10'd968: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller976;
		end
		10'd969: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller977;
		end
		10'd970: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller978;
		end
		10'd971: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller979;
		end
		10'd972: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller980;
		end
		10'd973: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller981;
		end
		10'd974: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller982;
		end
		10'd975: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller983;
		end
		10'd976: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller984;
		end
		10'd977: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller985;
		end
		10'd978: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller986;
		end
		10'd979: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller987;
		end
		10'd980: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller988;
		end
		10'd981: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller989;
		end
		10'd982: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller990;
		end
		10'd983: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller991;
		end
		10'd984: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller992;
		end
		10'd985: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller993;
		end
		10'd986: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller994;
		end
		10'd987: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller995;
		end
		10'd988: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller996;
		end
		10'd989: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller997;
		end
		10'd990: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller998;
		end
		10'd991: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller999;
		end
		10'd992: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1000;
		end
		10'd993: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1001;
		end
		10'd994: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1002;
		end
		10'd995: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1003;
		end
		10'd996: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1004;
		end
		10'd997: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1005;
		end
		10'd998: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1006;
		end
		10'd999: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1007;
		end
		10'd1000: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1008;
		end
		10'd1001: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1009;
		end
		10'd1002: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1010;
		end
		10'd1003: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1011;
		end
		10'd1004: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1012;
		end
		10'd1005: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1013;
		end
		10'd1006: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1014;
		end
		10'd1007: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1015;
		end
		10'd1008: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1016;
		end
		10'd1009: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1017;
		end
		10'd1010: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1018;
		end
		10'd1011: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1019;
		end
		10'd1012: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1020;
		end
		10'd1013: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1021;
		end
		10'd1014: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1022;
		end
		10'd1015: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1023;
		end
		10'd1016: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1024;
		end
		10'd1017: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1025;
		end
		10'd1018: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1026;
		end
		10'd1019: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1027;
		end
		10'd1020: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1028;
		end
		10'd1021: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1029;
		end
		10'd1022: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1030;
		end
		default: begin
			verilog_output_t_rhs_array_muxed <= mem_ctrl_memorycontroller1031;
		end
	endcase
// synthesis translate_off
	dummy_d_1 <= dummy_s;
// synthesis translate_on
end

// synthesis translate_off
reg dummy_d_2;
// synthesis translate_on
always @(*) begin
	verilog_output_f_rhs_array_muxed1 <= 64'd0;
	case (mem_ctrl_buffer_index)
		1'd0: begin
			verilog_output_f_rhs_array_muxed1 <= mem_ctrl_memorycontroller0;
		end
		1'd1: begin
			verilog_output_f_rhs_array_muxed1 <= mem_ctrl_memorycontroller1;
		end
		2'd2: begin
			verilog_output_f_rhs_array_muxed1 <= mem_ctrl_memorycontroller2;
		end
		2'd3: begin
			verilog_output_f_rhs_array_muxed1 <= mem_ctrl_memorycontroller3;
		end
		3'd4: begin
			verilog_output_f_rhs_array_muxed1 <= mem_ctrl_memorycontroller4;
		end
		3'd5: begin
			verilog_output_f_rhs_array_muxed1 <= mem_ctrl_memorycontroller5;
		end
		3'd6: begin
			verilog_output_f_rhs_array_muxed1 <= mem_ctrl_memorycontroller6;
		end
		default: begin
			verilog_output_f_rhs_array_muxed1 <= mem_ctrl_memorycontroller7;
		end
	endcase
// synthesis translate_off
	dummy_d_2 <= dummy_s;
// synthesis translate_on
end

always @(posedge sys_clk) begin
	if (rst) begin
		mem_ctrl_cmd_decoded <= 1'd0;
		mem_ctrl_address <= 1'd0;
	end else begin
		mem_ctrl_address <= addr;
		if (mem_read) begin
			mem_ctrl_cmd_decoded <= 2'd2;
		end else begin
			if (mem_write) begin
				mem_ctrl_cmd_decoded <= 2'd3;
			end else begin
				mem_ctrl_cmd_decoded <= 1'd0;
			end
		end
	end
	if (rst) begin
		mem_ctrl_timer <= 1'd0;
		mem_ctrl_state <= 1'd0;
		ready <= 1'd0;
	end else begin
		case (mem_ctrl_state)
			1'd0: begin
				if ((mem_ctrl_cmd_decoded != 1'd0)) begin
					mem_ctrl_state <= 1'd1;
					mem_ctrl_timer <= 1'd0;
					ready <= 1'd0;
				end
			end
			1'd1: begin
				if ((mem_ctrl_timer >= 4'd10)) begin
					mem_ctrl_state <= 2'd2;
					ready <= 1'd1;
				end else begin
					mem_ctrl_timer <= (mem_ctrl_timer + 1'd1);
				end
			end
			2'd2: begin
				mem_ctrl_state <= 1'd0;
			end
		endcase
	end
	if (rst) begin
		mem_ctrl_buffer_index <= 1'd0;
	end else begin
		if (ready) begin
			if (mem_write) begin
				verilog_output_t_lhs_array_muxed0 = data_in;
				case (mem_ctrl_buffer_index)
					1'd0: begin
						mem_ctrl_memorycontroller0 <= verilog_output_t_lhs_array_muxed0;
					end
					1'd1: begin
						mem_ctrl_memorycontroller1 <= verilog_output_t_lhs_array_muxed0;
					end
					2'd2: begin
						mem_ctrl_memorycontroller2 <= verilog_output_t_lhs_array_muxed0;
					end
					2'd3: begin
						mem_ctrl_memorycontroller3 <= verilog_output_t_lhs_array_muxed0;
					end
					3'd4: begin
						mem_ctrl_memorycontroller4 <= verilog_output_t_lhs_array_muxed0;
					end
					3'd5: begin
						mem_ctrl_memorycontroller5 <= verilog_output_t_lhs_array_muxed0;
					end
					3'd6: begin
						mem_ctrl_memorycontroller6 <= verilog_output_t_lhs_array_muxed0;
					end
					default: begin
						mem_ctrl_memorycontroller7 <= verilog_output_t_lhs_array_muxed0;
					end
				endcase
				if ((mem_ctrl_buffer_index == 3'd7)) begin
					mem_ctrl_buffer_index <= 1'd0;
				end else begin
					mem_ctrl_buffer_index <= (mem_ctrl_buffer_index + 1'd1);
				end
			end else begin
				if (mem_read) begin
					data_out <= verilog_output_f_rhs_array_muxed0;
					if ((mem_ctrl_buffer_index == 3'd7)) begin
						mem_ctrl_buffer_index <= 1'd0;
					end else begin
						mem_ctrl_buffer_index <= (mem_ctrl_buffer_index + 1'd1);
					end
				end
			end
		end
	end
	if (rst) begin
		mem_ctrl_power_state <= 1'd0;
	end else begin
		case (mem_ctrl_power_state)
			1'd0: begin
				if ((mem_ctrl_cmd_decoded == 1'd0)) begin
					mem_ctrl_power_state <= 1'd1;
				end
			end
			1'd1: begin
				if ((mem_ctrl_cmd_decoded != 1'd0)) begin
					mem_ctrl_power_state <= 1'd0;
				end
			end
		endcase
	end
	if (rst) begin
	end else begin
		if (ready) begin
			if (mem_read) begin
				verilog_output_t_lhs_array_muxed1 = verilog_output_t_rhs_array_muxed;
				case (mem_ctrl_buffer_index)
					1'd0: begin
						mem_ctrl_memorycontroller0 <= verilog_output_t_lhs_array_muxed1;
					end
					1'd1: begin
						mem_ctrl_memorycontroller1 <= verilog_output_t_lhs_array_muxed1;
					end
					2'd2: begin
						mem_ctrl_memorycontroller2 <= verilog_output_t_lhs_array_muxed1;
					end
					2'd3: begin
						mem_ctrl_memorycontroller3 <= verilog_output_t_lhs_array_muxed1;
					end
					3'd4: begin
						mem_ctrl_memorycontroller4 <= verilog_output_t_lhs_array_muxed1;
					end
					3'd5: begin
						mem_ctrl_memorycontroller5 <= verilog_output_t_lhs_array_muxed1;
					end
					3'd6: begin
						mem_ctrl_memorycontroller6 <= verilog_output_t_lhs_array_muxed1;
					end
					default: begin
						mem_ctrl_memorycontroller7 <= verilog_output_t_lhs_array_muxed1;
					end
				endcase
			end else begin
				if (mem_write) begin
					verilog_output_f_lhs_array_muxed = verilog_output_f_rhs_array_muxed1;
					case (mem_ctrl_address)
						1'd0: begin
							mem_ctrl_memorycontroller8 <= verilog_output_f_lhs_array_muxed;
						end
						1'd1: begin
							mem_ctrl_memorycontroller9 <= verilog_output_f_lhs_array_muxed;
						end
						2'd2: begin
							mem_ctrl_memorycontroller10 <= verilog_output_f_lhs_array_muxed;
						end
						2'd3: begin
							mem_ctrl_memorycontroller11 <= verilog_output_f_lhs_array_muxed;
						end
						3'd4: begin
							mem_ctrl_memorycontroller12 <= verilog_output_f_lhs_array_muxed;
						end
						3'd5: begin
							mem_ctrl_memorycontroller13 <= verilog_output_f_lhs_array_muxed;
						end
						3'd6: begin
							mem_ctrl_memorycontroller14 <= verilog_output_f_lhs_array_muxed;
						end
						3'd7: begin
							mem_ctrl_memorycontroller15 <= verilog_output_f_lhs_array_muxed;
						end
						4'd8: begin
							mem_ctrl_memorycontroller16 <= verilog_output_f_lhs_array_muxed;
						end
						4'd9: begin
							mem_ctrl_memorycontroller17 <= verilog_output_f_lhs_array_muxed;
						end
						4'd10: begin
							mem_ctrl_memorycontroller18 <= verilog_output_f_lhs_array_muxed;
						end
						4'd11: begin
							mem_ctrl_memorycontroller19 <= verilog_output_f_lhs_array_muxed;
						end
						4'd12: begin
							mem_ctrl_memorycontroller20 <= verilog_output_f_lhs_array_muxed;
						end
						4'd13: begin
							mem_ctrl_memorycontroller21 <= verilog_output_f_lhs_array_muxed;
						end
						4'd14: begin
							mem_ctrl_memorycontroller22 <= verilog_output_f_lhs_array_muxed;
						end
						4'd15: begin
							mem_ctrl_memorycontroller23 <= verilog_output_f_lhs_array_muxed;
						end
						5'd16: begin
							mem_ctrl_memorycontroller24 <= verilog_output_f_lhs_array_muxed;
						end
						5'd17: begin
							mem_ctrl_memorycontroller25 <= verilog_output_f_lhs_array_muxed;
						end
						5'd18: begin
							mem_ctrl_memorycontroller26 <= verilog_output_f_lhs_array_muxed;
						end
						5'd19: begin
							mem_ctrl_memorycontroller27 <= verilog_output_f_lhs_array_muxed;
						end
						5'd20: begin
							mem_ctrl_memorycontroller28 <= verilog_output_f_lhs_array_muxed;
						end
						5'd21: begin
							mem_ctrl_memorycontroller29 <= verilog_output_f_lhs_array_muxed;
						end
						5'd22: begin
							mem_ctrl_memorycontroller30 <= verilog_output_f_lhs_array_muxed;
						end
						5'd23: begin
							mem_ctrl_memorycontroller31 <= verilog_output_f_lhs_array_muxed;
						end
						5'd24: begin
							mem_ctrl_memorycontroller32 <= verilog_output_f_lhs_array_muxed;
						end
						5'd25: begin
							mem_ctrl_memorycontroller33 <= verilog_output_f_lhs_array_muxed;
						end
						5'd26: begin
							mem_ctrl_memorycontroller34 <= verilog_output_f_lhs_array_muxed;
						end
						5'd27: begin
							mem_ctrl_memorycontroller35 <= verilog_output_f_lhs_array_muxed;
						end
						5'd28: begin
							mem_ctrl_memorycontroller36 <= verilog_output_f_lhs_array_muxed;
						end
						5'd29: begin
							mem_ctrl_memorycontroller37 <= verilog_output_f_lhs_array_muxed;
						end
						5'd30: begin
							mem_ctrl_memorycontroller38 <= verilog_output_f_lhs_array_muxed;
						end
						5'd31: begin
							mem_ctrl_memorycontroller39 <= verilog_output_f_lhs_array_muxed;
						end
						6'd32: begin
							mem_ctrl_memorycontroller40 <= verilog_output_f_lhs_array_muxed;
						end
						6'd33: begin
							mem_ctrl_memorycontroller41 <= verilog_output_f_lhs_array_muxed;
						end
						6'd34: begin
							mem_ctrl_memorycontroller42 <= verilog_output_f_lhs_array_muxed;
						end
						6'd35: begin
							mem_ctrl_memorycontroller43 <= verilog_output_f_lhs_array_muxed;
						end
						6'd36: begin
							mem_ctrl_memorycontroller44 <= verilog_output_f_lhs_array_muxed;
						end
						6'd37: begin
							mem_ctrl_memorycontroller45 <= verilog_output_f_lhs_array_muxed;
						end
						6'd38: begin
							mem_ctrl_memorycontroller46 <= verilog_output_f_lhs_array_muxed;
						end
						6'd39: begin
							mem_ctrl_memorycontroller47 <= verilog_output_f_lhs_array_muxed;
						end
						6'd40: begin
							mem_ctrl_memorycontroller48 <= verilog_output_f_lhs_array_muxed;
						end
						6'd41: begin
							mem_ctrl_memorycontroller49 <= verilog_output_f_lhs_array_muxed;
						end
						6'd42: begin
							mem_ctrl_memorycontroller50 <= verilog_output_f_lhs_array_muxed;
						end
						6'd43: begin
							mem_ctrl_memorycontroller51 <= verilog_output_f_lhs_array_muxed;
						end
						6'd44: begin
							mem_ctrl_memorycontroller52 <= verilog_output_f_lhs_array_muxed;
						end
						6'd45: begin
							mem_ctrl_memorycontroller53 <= verilog_output_f_lhs_array_muxed;
						end
						6'd46: begin
							mem_ctrl_memorycontroller54 <= verilog_output_f_lhs_array_muxed;
						end
						6'd47: begin
							mem_ctrl_memorycontroller55 <= verilog_output_f_lhs_array_muxed;
						end
						6'd48: begin
							mem_ctrl_memorycontroller56 <= verilog_output_f_lhs_array_muxed;
						end
						6'd49: begin
							mem_ctrl_memorycontroller57 <= verilog_output_f_lhs_array_muxed;
						end
						6'd50: begin
							mem_ctrl_memorycontroller58 <= verilog_output_f_lhs_array_muxed;
						end
						6'd51: begin
							mem_ctrl_memorycontroller59 <= verilog_output_f_lhs_array_muxed;
						end
						6'd52: begin
							mem_ctrl_memorycontroller60 <= verilog_output_f_lhs_array_muxed;
						end
						6'd53: begin
							mem_ctrl_memorycontroller61 <= verilog_output_f_lhs_array_muxed;
						end
						6'd54: begin
							mem_ctrl_memorycontroller62 <= verilog_output_f_lhs_array_muxed;
						end
						6'd55: begin
							mem_ctrl_memorycontroller63 <= verilog_output_f_lhs_array_muxed;
						end
						6'd56: begin
							mem_ctrl_memorycontroller64 <= verilog_output_f_lhs_array_muxed;
						end
						6'd57: begin
							mem_ctrl_memorycontroller65 <= verilog_output_f_lhs_array_muxed;
						end
						6'd58: begin
							mem_ctrl_memorycontroller66 <= verilog_output_f_lhs_array_muxed;
						end
						6'd59: begin
							mem_ctrl_memorycontroller67 <= verilog_output_f_lhs_array_muxed;
						end
						6'd60: begin
							mem_ctrl_memorycontroller68 <= verilog_output_f_lhs_array_muxed;
						end
						6'd61: begin
							mem_ctrl_memorycontroller69 <= verilog_output_f_lhs_array_muxed;
						end
						6'd62: begin
							mem_ctrl_memorycontroller70 <= verilog_output_f_lhs_array_muxed;
						end
						6'd63: begin
							mem_ctrl_memorycontroller71 <= verilog_output_f_lhs_array_muxed;
						end
						7'd64: begin
							mem_ctrl_memorycontroller72 <= verilog_output_f_lhs_array_muxed;
						end
						7'd65: begin
							mem_ctrl_memorycontroller73 <= verilog_output_f_lhs_array_muxed;
						end
						7'd66: begin
							mem_ctrl_memorycontroller74 <= verilog_output_f_lhs_array_muxed;
						end
						7'd67: begin
							mem_ctrl_memorycontroller75 <= verilog_output_f_lhs_array_muxed;
						end
						7'd68: begin
							mem_ctrl_memorycontroller76 <= verilog_output_f_lhs_array_muxed;
						end
						7'd69: begin
							mem_ctrl_memorycontroller77 <= verilog_output_f_lhs_array_muxed;
						end
						7'd70: begin
							mem_ctrl_memorycontroller78 <= verilog_output_f_lhs_array_muxed;
						end
						7'd71: begin
							mem_ctrl_memorycontroller79 <= verilog_output_f_lhs_array_muxed;
						end
						7'd72: begin
							mem_ctrl_memorycontroller80 <= verilog_output_f_lhs_array_muxed;
						end
						7'd73: begin
							mem_ctrl_memorycontroller81 <= verilog_output_f_lhs_array_muxed;
						end
						7'd74: begin
							mem_ctrl_memorycontroller82 <= verilog_output_f_lhs_array_muxed;
						end
						7'd75: begin
							mem_ctrl_memorycontroller83 <= verilog_output_f_lhs_array_muxed;
						end
						7'd76: begin
							mem_ctrl_memorycontroller84 <= verilog_output_f_lhs_array_muxed;
						end
						7'd77: begin
							mem_ctrl_memorycontroller85 <= verilog_output_f_lhs_array_muxed;
						end
						7'd78: begin
							mem_ctrl_memorycontroller86 <= verilog_output_f_lhs_array_muxed;
						end
						7'd79: begin
							mem_ctrl_memorycontroller87 <= verilog_output_f_lhs_array_muxed;
						end
						7'd80: begin
							mem_ctrl_memorycontroller88 <= verilog_output_f_lhs_array_muxed;
						end
						7'd81: begin
							mem_ctrl_memorycontroller89 <= verilog_output_f_lhs_array_muxed;
						end
						7'd82: begin
							mem_ctrl_memorycontroller90 <= verilog_output_f_lhs_array_muxed;
						end
						7'd83: begin
							mem_ctrl_memorycontroller91 <= verilog_output_f_lhs_array_muxed;
						end
						7'd84: begin
							mem_ctrl_memorycontroller92 <= verilog_output_f_lhs_array_muxed;
						end
						7'd85: begin
							mem_ctrl_memorycontroller93 <= verilog_output_f_lhs_array_muxed;
						end
						7'd86: begin
							mem_ctrl_memorycontroller94 <= verilog_output_f_lhs_array_muxed;
						end
						7'd87: begin
							mem_ctrl_memorycontroller95 <= verilog_output_f_lhs_array_muxed;
						end
						7'd88: begin
							mem_ctrl_memorycontroller96 <= verilog_output_f_lhs_array_muxed;
						end
						7'd89: begin
							mem_ctrl_memorycontroller97 <= verilog_output_f_lhs_array_muxed;
						end
						7'd90: begin
							mem_ctrl_memorycontroller98 <= verilog_output_f_lhs_array_muxed;
						end
						7'd91: begin
							mem_ctrl_memorycontroller99 <= verilog_output_f_lhs_array_muxed;
						end
						7'd92: begin
							mem_ctrl_memorycontroller100 <= verilog_output_f_lhs_array_muxed;
						end
						7'd93: begin
							mem_ctrl_memorycontroller101 <= verilog_output_f_lhs_array_muxed;
						end
						7'd94: begin
							mem_ctrl_memorycontroller102 <= verilog_output_f_lhs_array_muxed;
						end
						7'd95: begin
							mem_ctrl_memorycontroller103 <= verilog_output_f_lhs_array_muxed;
						end
						7'd96: begin
							mem_ctrl_memorycontroller104 <= verilog_output_f_lhs_array_muxed;
						end
						7'd97: begin
							mem_ctrl_memorycontroller105 <= verilog_output_f_lhs_array_muxed;
						end
						7'd98: begin
							mem_ctrl_memorycontroller106 <= verilog_output_f_lhs_array_muxed;
						end
						7'd99: begin
							mem_ctrl_memorycontroller107 <= verilog_output_f_lhs_array_muxed;
						end
						7'd100: begin
							mem_ctrl_memorycontroller108 <= verilog_output_f_lhs_array_muxed;
						end
						7'd101: begin
							mem_ctrl_memorycontroller109 <= verilog_output_f_lhs_array_muxed;
						end
						7'd102: begin
							mem_ctrl_memorycontroller110 <= verilog_output_f_lhs_array_muxed;
						end
						7'd103: begin
							mem_ctrl_memorycontroller111 <= verilog_output_f_lhs_array_muxed;
						end
						7'd104: begin
							mem_ctrl_memorycontroller112 <= verilog_output_f_lhs_array_muxed;
						end
						7'd105: begin
							mem_ctrl_memorycontroller113 <= verilog_output_f_lhs_array_muxed;
						end
						7'd106: begin
							mem_ctrl_memorycontroller114 <= verilog_output_f_lhs_array_muxed;
						end
						7'd107: begin
							mem_ctrl_memorycontroller115 <= verilog_output_f_lhs_array_muxed;
						end
						7'd108: begin
							mem_ctrl_memorycontroller116 <= verilog_output_f_lhs_array_muxed;
						end
						7'd109: begin
							mem_ctrl_memorycontroller117 <= verilog_output_f_lhs_array_muxed;
						end
						7'd110: begin
							mem_ctrl_memorycontroller118 <= verilog_output_f_lhs_array_muxed;
						end
						7'd111: begin
							mem_ctrl_memorycontroller119 <= verilog_output_f_lhs_array_muxed;
						end
						7'd112: begin
							mem_ctrl_memorycontroller120 <= verilog_output_f_lhs_array_muxed;
						end
						7'd113: begin
							mem_ctrl_memorycontroller121 <= verilog_output_f_lhs_array_muxed;
						end
						7'd114: begin
							mem_ctrl_memorycontroller122 <= verilog_output_f_lhs_array_muxed;
						end
						7'd115: begin
							mem_ctrl_memorycontroller123 <= verilog_output_f_lhs_array_muxed;
						end
						7'd116: begin
							mem_ctrl_memorycontroller124 <= verilog_output_f_lhs_array_muxed;
						end
						7'd117: begin
							mem_ctrl_memorycontroller125 <= verilog_output_f_lhs_array_muxed;
						end
						7'd118: begin
							mem_ctrl_memorycontroller126 <= verilog_output_f_lhs_array_muxed;
						end
						7'd119: begin
							mem_ctrl_memorycontroller127 <= verilog_output_f_lhs_array_muxed;
						end
						7'd120: begin
							mem_ctrl_memorycontroller128 <= verilog_output_f_lhs_array_muxed;
						end
						7'd121: begin
							mem_ctrl_memorycontroller129 <= verilog_output_f_lhs_array_muxed;
						end
						7'd122: begin
							mem_ctrl_memorycontroller130 <= verilog_output_f_lhs_array_muxed;
						end
						7'd123: begin
							mem_ctrl_memorycontroller131 <= verilog_output_f_lhs_array_muxed;
						end
						7'd124: begin
							mem_ctrl_memorycontroller132 <= verilog_output_f_lhs_array_muxed;
						end
						7'd125: begin
							mem_ctrl_memorycontroller133 <= verilog_output_f_lhs_array_muxed;
						end
						7'd126: begin
							mem_ctrl_memorycontroller134 <= verilog_output_f_lhs_array_muxed;
						end
						7'd127: begin
							mem_ctrl_memorycontroller135 <= verilog_output_f_lhs_array_muxed;
						end
						8'd128: begin
							mem_ctrl_memorycontroller136 <= verilog_output_f_lhs_array_muxed;
						end
						8'd129: begin
							mem_ctrl_memorycontroller137 <= verilog_output_f_lhs_array_muxed;
						end
						8'd130: begin
							mem_ctrl_memorycontroller138 <= verilog_output_f_lhs_array_muxed;
						end
						8'd131: begin
							mem_ctrl_memorycontroller139 <= verilog_output_f_lhs_array_muxed;
						end
						8'd132: begin
							mem_ctrl_memorycontroller140 <= verilog_output_f_lhs_array_muxed;
						end
						8'd133: begin
							mem_ctrl_memorycontroller141 <= verilog_output_f_lhs_array_muxed;
						end
						8'd134: begin
							mem_ctrl_memorycontroller142 <= verilog_output_f_lhs_array_muxed;
						end
						8'd135: begin
							mem_ctrl_memorycontroller143 <= verilog_output_f_lhs_array_muxed;
						end
						8'd136: begin
							mem_ctrl_memorycontroller144 <= verilog_output_f_lhs_array_muxed;
						end
						8'd137: begin
							mem_ctrl_memorycontroller145 <= verilog_output_f_lhs_array_muxed;
						end
						8'd138: begin
							mem_ctrl_memorycontroller146 <= verilog_output_f_lhs_array_muxed;
						end
						8'd139: begin
							mem_ctrl_memorycontroller147 <= verilog_output_f_lhs_array_muxed;
						end
						8'd140: begin
							mem_ctrl_memorycontroller148 <= verilog_output_f_lhs_array_muxed;
						end
						8'd141: begin
							mem_ctrl_memorycontroller149 <= verilog_output_f_lhs_array_muxed;
						end
						8'd142: begin
							mem_ctrl_memorycontroller150 <= verilog_output_f_lhs_array_muxed;
						end
						8'd143: begin
							mem_ctrl_memorycontroller151 <= verilog_output_f_lhs_array_muxed;
						end
						8'd144: begin
							mem_ctrl_memorycontroller152 <= verilog_output_f_lhs_array_muxed;
						end
						8'd145: begin
							mem_ctrl_memorycontroller153 <= verilog_output_f_lhs_array_muxed;
						end
						8'd146: begin
							mem_ctrl_memorycontroller154 <= verilog_output_f_lhs_array_muxed;
						end
						8'd147: begin
							mem_ctrl_memorycontroller155 <= verilog_output_f_lhs_array_muxed;
						end
						8'd148: begin
							mem_ctrl_memorycontroller156 <= verilog_output_f_lhs_array_muxed;
						end
						8'd149: begin
							mem_ctrl_memorycontroller157 <= verilog_output_f_lhs_array_muxed;
						end
						8'd150: begin
							mem_ctrl_memorycontroller158 <= verilog_output_f_lhs_array_muxed;
						end
						8'd151: begin
							mem_ctrl_memorycontroller159 <= verilog_output_f_lhs_array_muxed;
						end
						8'd152: begin
							mem_ctrl_memorycontroller160 <= verilog_output_f_lhs_array_muxed;
						end
						8'd153: begin
							mem_ctrl_memorycontroller161 <= verilog_output_f_lhs_array_muxed;
						end
						8'd154: begin
							mem_ctrl_memorycontroller162 <= verilog_output_f_lhs_array_muxed;
						end
						8'd155: begin
							mem_ctrl_memorycontroller163 <= verilog_output_f_lhs_array_muxed;
						end
						8'd156: begin
							mem_ctrl_memorycontroller164 <= verilog_output_f_lhs_array_muxed;
						end
						8'd157: begin
							mem_ctrl_memorycontroller165 <= verilog_output_f_lhs_array_muxed;
						end
						8'd158: begin
							mem_ctrl_memorycontroller166 <= verilog_output_f_lhs_array_muxed;
						end
						8'd159: begin
							mem_ctrl_memorycontroller167 <= verilog_output_f_lhs_array_muxed;
						end
						8'd160: begin
							mem_ctrl_memorycontroller168 <= verilog_output_f_lhs_array_muxed;
						end
						8'd161: begin
							mem_ctrl_memorycontroller169 <= verilog_output_f_lhs_array_muxed;
						end
						8'd162: begin
							mem_ctrl_memorycontroller170 <= verilog_output_f_lhs_array_muxed;
						end
						8'd163: begin
							mem_ctrl_memorycontroller171 <= verilog_output_f_lhs_array_muxed;
						end
						8'd164: begin
							mem_ctrl_memorycontroller172 <= verilog_output_f_lhs_array_muxed;
						end
						8'd165: begin
							mem_ctrl_memorycontroller173 <= verilog_output_f_lhs_array_muxed;
						end
						8'd166: begin
							mem_ctrl_memorycontroller174 <= verilog_output_f_lhs_array_muxed;
						end
						8'd167: begin
							mem_ctrl_memorycontroller175 <= verilog_output_f_lhs_array_muxed;
						end
						8'd168: begin
							mem_ctrl_memorycontroller176 <= verilog_output_f_lhs_array_muxed;
						end
						8'd169: begin
							mem_ctrl_memorycontroller177 <= verilog_output_f_lhs_array_muxed;
						end
						8'd170: begin
							mem_ctrl_memorycontroller178 <= verilog_output_f_lhs_array_muxed;
						end
						8'd171: begin
							mem_ctrl_memorycontroller179 <= verilog_output_f_lhs_array_muxed;
						end
						8'd172: begin
							mem_ctrl_memorycontroller180 <= verilog_output_f_lhs_array_muxed;
						end
						8'd173: begin
							mem_ctrl_memorycontroller181 <= verilog_output_f_lhs_array_muxed;
						end
						8'd174: begin
							mem_ctrl_memorycontroller182 <= verilog_output_f_lhs_array_muxed;
						end
						8'd175: begin
							mem_ctrl_memorycontroller183 <= verilog_output_f_lhs_array_muxed;
						end
						8'd176: begin
							mem_ctrl_memorycontroller184 <= verilog_output_f_lhs_array_muxed;
						end
						8'd177: begin
							mem_ctrl_memorycontroller185 <= verilog_output_f_lhs_array_muxed;
						end
						8'd178: begin
							mem_ctrl_memorycontroller186 <= verilog_output_f_lhs_array_muxed;
						end
						8'd179: begin
							mem_ctrl_memorycontroller187 <= verilog_output_f_lhs_array_muxed;
						end
						8'd180: begin
							mem_ctrl_memorycontroller188 <= verilog_output_f_lhs_array_muxed;
						end
						8'd181: begin
							mem_ctrl_memorycontroller189 <= verilog_output_f_lhs_array_muxed;
						end
						8'd182: begin
							mem_ctrl_memorycontroller190 <= verilog_output_f_lhs_array_muxed;
						end
						8'd183: begin
							mem_ctrl_memorycontroller191 <= verilog_output_f_lhs_array_muxed;
						end
						8'd184: begin
							mem_ctrl_memorycontroller192 <= verilog_output_f_lhs_array_muxed;
						end
						8'd185: begin
							mem_ctrl_memorycontroller193 <= verilog_output_f_lhs_array_muxed;
						end
						8'd186: begin
							mem_ctrl_memorycontroller194 <= verilog_output_f_lhs_array_muxed;
						end
						8'd187: begin
							mem_ctrl_memorycontroller195 <= verilog_output_f_lhs_array_muxed;
						end
						8'd188: begin
							mem_ctrl_memorycontroller196 <= verilog_output_f_lhs_array_muxed;
						end
						8'd189: begin
							mem_ctrl_memorycontroller197 <= verilog_output_f_lhs_array_muxed;
						end
						8'd190: begin
							mem_ctrl_memorycontroller198 <= verilog_output_f_lhs_array_muxed;
						end
						8'd191: begin
							mem_ctrl_memorycontroller199 <= verilog_output_f_lhs_array_muxed;
						end
						8'd192: begin
							mem_ctrl_memorycontroller200 <= verilog_output_f_lhs_array_muxed;
						end
						8'd193: begin
							mem_ctrl_memorycontroller201 <= verilog_output_f_lhs_array_muxed;
						end
						8'd194: begin
							mem_ctrl_memorycontroller202 <= verilog_output_f_lhs_array_muxed;
						end
						8'd195: begin
							mem_ctrl_memorycontroller203 <= verilog_output_f_lhs_array_muxed;
						end
						8'd196: begin
							mem_ctrl_memorycontroller204 <= verilog_output_f_lhs_array_muxed;
						end
						8'd197: begin
							mem_ctrl_memorycontroller205 <= verilog_output_f_lhs_array_muxed;
						end
						8'd198: begin
							mem_ctrl_memorycontroller206 <= verilog_output_f_lhs_array_muxed;
						end
						8'd199: begin
							mem_ctrl_memorycontroller207 <= verilog_output_f_lhs_array_muxed;
						end
						8'd200: begin
							mem_ctrl_memorycontroller208 <= verilog_output_f_lhs_array_muxed;
						end
						8'd201: begin
							mem_ctrl_memorycontroller209 <= verilog_output_f_lhs_array_muxed;
						end
						8'd202: begin
							mem_ctrl_memorycontroller210 <= verilog_output_f_lhs_array_muxed;
						end
						8'd203: begin
							mem_ctrl_memorycontroller211 <= verilog_output_f_lhs_array_muxed;
						end
						8'd204: begin
							mem_ctrl_memorycontroller212 <= verilog_output_f_lhs_array_muxed;
						end
						8'd205: begin
							mem_ctrl_memorycontroller213 <= verilog_output_f_lhs_array_muxed;
						end
						8'd206: begin
							mem_ctrl_memorycontroller214 <= verilog_output_f_lhs_array_muxed;
						end
						8'd207: begin
							mem_ctrl_memorycontroller215 <= verilog_output_f_lhs_array_muxed;
						end
						8'd208: begin
							mem_ctrl_memorycontroller216 <= verilog_output_f_lhs_array_muxed;
						end
						8'd209: begin
							mem_ctrl_memorycontroller217 <= verilog_output_f_lhs_array_muxed;
						end
						8'd210: begin
							mem_ctrl_memorycontroller218 <= verilog_output_f_lhs_array_muxed;
						end
						8'd211: begin
							mem_ctrl_memorycontroller219 <= verilog_output_f_lhs_array_muxed;
						end
						8'd212: begin
							mem_ctrl_memorycontroller220 <= verilog_output_f_lhs_array_muxed;
						end
						8'd213: begin
							mem_ctrl_memorycontroller221 <= verilog_output_f_lhs_array_muxed;
						end
						8'd214: begin
							mem_ctrl_memorycontroller222 <= verilog_output_f_lhs_array_muxed;
						end
						8'd215: begin
							mem_ctrl_memorycontroller223 <= verilog_output_f_lhs_array_muxed;
						end
						8'd216: begin
							mem_ctrl_memorycontroller224 <= verilog_output_f_lhs_array_muxed;
						end
						8'd217: begin
							mem_ctrl_memorycontroller225 <= verilog_output_f_lhs_array_muxed;
						end
						8'd218: begin
							mem_ctrl_memorycontroller226 <= verilog_output_f_lhs_array_muxed;
						end
						8'd219: begin
							mem_ctrl_memorycontroller227 <= verilog_output_f_lhs_array_muxed;
						end
						8'd220: begin
							mem_ctrl_memorycontroller228 <= verilog_output_f_lhs_array_muxed;
						end
						8'd221: begin
							mem_ctrl_memorycontroller229 <= verilog_output_f_lhs_array_muxed;
						end
						8'd222: begin
							mem_ctrl_memorycontroller230 <= verilog_output_f_lhs_array_muxed;
						end
						8'd223: begin
							mem_ctrl_memorycontroller231 <= verilog_output_f_lhs_array_muxed;
						end
						8'd224: begin
							mem_ctrl_memorycontroller232 <= verilog_output_f_lhs_array_muxed;
						end
						8'd225: begin
							mem_ctrl_memorycontroller233 <= verilog_output_f_lhs_array_muxed;
						end
						8'd226: begin
							mem_ctrl_memorycontroller234 <= verilog_output_f_lhs_array_muxed;
						end
						8'd227: begin
							mem_ctrl_memorycontroller235 <= verilog_output_f_lhs_array_muxed;
						end
						8'd228: begin
							mem_ctrl_memorycontroller236 <= verilog_output_f_lhs_array_muxed;
						end
						8'd229: begin
							mem_ctrl_memorycontroller237 <= verilog_output_f_lhs_array_muxed;
						end
						8'd230: begin
							mem_ctrl_memorycontroller238 <= verilog_output_f_lhs_array_muxed;
						end
						8'd231: begin
							mem_ctrl_memorycontroller239 <= verilog_output_f_lhs_array_muxed;
						end
						8'd232: begin
							mem_ctrl_memorycontroller240 <= verilog_output_f_lhs_array_muxed;
						end
						8'd233: begin
							mem_ctrl_memorycontroller241 <= verilog_output_f_lhs_array_muxed;
						end
						8'd234: begin
							mem_ctrl_memorycontroller242 <= verilog_output_f_lhs_array_muxed;
						end
						8'd235: begin
							mem_ctrl_memorycontroller243 <= verilog_output_f_lhs_array_muxed;
						end
						8'd236: begin
							mem_ctrl_memorycontroller244 <= verilog_output_f_lhs_array_muxed;
						end
						8'd237: begin
							mem_ctrl_memorycontroller245 <= verilog_output_f_lhs_array_muxed;
						end
						8'd238: begin
							mem_ctrl_memorycontroller246 <= verilog_output_f_lhs_array_muxed;
						end
						8'd239: begin
							mem_ctrl_memorycontroller247 <= verilog_output_f_lhs_array_muxed;
						end
						8'd240: begin
							mem_ctrl_memorycontroller248 <= verilog_output_f_lhs_array_muxed;
						end
						8'd241: begin
							mem_ctrl_memorycontroller249 <= verilog_output_f_lhs_array_muxed;
						end
						8'd242: begin
							mem_ctrl_memorycontroller250 <= verilog_output_f_lhs_array_muxed;
						end
						8'd243: begin
							mem_ctrl_memorycontroller251 <= verilog_output_f_lhs_array_muxed;
						end
						8'd244: begin
							mem_ctrl_memorycontroller252 <= verilog_output_f_lhs_array_muxed;
						end
						8'd245: begin
							mem_ctrl_memorycontroller253 <= verilog_output_f_lhs_array_muxed;
						end
						8'd246: begin
							mem_ctrl_memorycontroller254 <= verilog_output_f_lhs_array_muxed;
						end
						8'd247: begin
							mem_ctrl_memorycontroller255 <= verilog_output_f_lhs_array_muxed;
						end
						8'd248: begin
							mem_ctrl_memorycontroller256 <= verilog_output_f_lhs_array_muxed;
						end
						8'd249: begin
							mem_ctrl_memorycontroller257 <= verilog_output_f_lhs_array_muxed;
						end
						8'd250: begin
							mem_ctrl_memorycontroller258 <= verilog_output_f_lhs_array_muxed;
						end
						8'd251: begin
							mem_ctrl_memorycontroller259 <= verilog_output_f_lhs_array_muxed;
						end
						8'd252: begin
							mem_ctrl_memorycontroller260 <= verilog_output_f_lhs_array_muxed;
						end
						8'd253: begin
							mem_ctrl_memorycontroller261 <= verilog_output_f_lhs_array_muxed;
						end
						8'd254: begin
							mem_ctrl_memorycontroller262 <= verilog_output_f_lhs_array_muxed;
						end
						8'd255: begin
							mem_ctrl_memorycontroller263 <= verilog_output_f_lhs_array_muxed;
						end
						9'd256: begin
							mem_ctrl_memorycontroller264 <= verilog_output_f_lhs_array_muxed;
						end
						9'd257: begin
							mem_ctrl_memorycontroller265 <= verilog_output_f_lhs_array_muxed;
						end
						9'd258: begin
							mem_ctrl_memorycontroller266 <= verilog_output_f_lhs_array_muxed;
						end
						9'd259: begin
							mem_ctrl_memorycontroller267 <= verilog_output_f_lhs_array_muxed;
						end
						9'd260: begin
							mem_ctrl_memorycontroller268 <= verilog_output_f_lhs_array_muxed;
						end
						9'd261: begin
							mem_ctrl_memorycontroller269 <= verilog_output_f_lhs_array_muxed;
						end
						9'd262: begin
							mem_ctrl_memorycontroller270 <= verilog_output_f_lhs_array_muxed;
						end
						9'd263: begin
							mem_ctrl_memorycontroller271 <= verilog_output_f_lhs_array_muxed;
						end
						9'd264: begin
							mem_ctrl_memorycontroller272 <= verilog_output_f_lhs_array_muxed;
						end
						9'd265: begin
							mem_ctrl_memorycontroller273 <= verilog_output_f_lhs_array_muxed;
						end
						9'd266: begin
							mem_ctrl_memorycontroller274 <= verilog_output_f_lhs_array_muxed;
						end
						9'd267: begin
							mem_ctrl_memorycontroller275 <= verilog_output_f_lhs_array_muxed;
						end
						9'd268: begin
							mem_ctrl_memorycontroller276 <= verilog_output_f_lhs_array_muxed;
						end
						9'd269: begin
							mem_ctrl_memorycontroller277 <= verilog_output_f_lhs_array_muxed;
						end
						9'd270: begin
							mem_ctrl_memorycontroller278 <= verilog_output_f_lhs_array_muxed;
						end
						9'd271: begin
							mem_ctrl_memorycontroller279 <= verilog_output_f_lhs_array_muxed;
						end
						9'd272: begin
							mem_ctrl_memorycontroller280 <= verilog_output_f_lhs_array_muxed;
						end
						9'd273: begin
							mem_ctrl_memorycontroller281 <= verilog_output_f_lhs_array_muxed;
						end
						9'd274: begin
							mem_ctrl_memorycontroller282 <= verilog_output_f_lhs_array_muxed;
						end
						9'd275: begin
							mem_ctrl_memorycontroller283 <= verilog_output_f_lhs_array_muxed;
						end
						9'd276: begin
							mem_ctrl_memorycontroller284 <= verilog_output_f_lhs_array_muxed;
						end
						9'd277: begin
							mem_ctrl_memorycontroller285 <= verilog_output_f_lhs_array_muxed;
						end
						9'd278: begin
							mem_ctrl_memorycontroller286 <= verilog_output_f_lhs_array_muxed;
						end
						9'd279: begin
							mem_ctrl_memorycontroller287 <= verilog_output_f_lhs_array_muxed;
						end
						9'd280: begin
							mem_ctrl_memorycontroller288 <= verilog_output_f_lhs_array_muxed;
						end
						9'd281: begin
							mem_ctrl_memorycontroller289 <= verilog_output_f_lhs_array_muxed;
						end
						9'd282: begin
							mem_ctrl_memorycontroller290 <= verilog_output_f_lhs_array_muxed;
						end
						9'd283: begin
							mem_ctrl_memorycontroller291 <= verilog_output_f_lhs_array_muxed;
						end
						9'd284: begin
							mem_ctrl_memorycontroller292 <= verilog_output_f_lhs_array_muxed;
						end
						9'd285: begin
							mem_ctrl_memorycontroller293 <= verilog_output_f_lhs_array_muxed;
						end
						9'd286: begin
							mem_ctrl_memorycontroller294 <= verilog_output_f_lhs_array_muxed;
						end
						9'd287: begin
							mem_ctrl_memorycontroller295 <= verilog_output_f_lhs_array_muxed;
						end
						9'd288: begin
							mem_ctrl_memorycontroller296 <= verilog_output_f_lhs_array_muxed;
						end
						9'd289: begin
							mem_ctrl_memorycontroller297 <= verilog_output_f_lhs_array_muxed;
						end
						9'd290: begin
							mem_ctrl_memorycontroller298 <= verilog_output_f_lhs_array_muxed;
						end
						9'd291: begin
							mem_ctrl_memorycontroller299 <= verilog_output_f_lhs_array_muxed;
						end
						9'd292: begin
							mem_ctrl_memorycontroller300 <= verilog_output_f_lhs_array_muxed;
						end
						9'd293: begin
							mem_ctrl_memorycontroller301 <= verilog_output_f_lhs_array_muxed;
						end
						9'd294: begin
							mem_ctrl_memorycontroller302 <= verilog_output_f_lhs_array_muxed;
						end
						9'd295: begin
							mem_ctrl_memorycontroller303 <= verilog_output_f_lhs_array_muxed;
						end
						9'd296: begin
							mem_ctrl_memorycontroller304 <= verilog_output_f_lhs_array_muxed;
						end
						9'd297: begin
							mem_ctrl_memorycontroller305 <= verilog_output_f_lhs_array_muxed;
						end
						9'd298: begin
							mem_ctrl_memorycontroller306 <= verilog_output_f_lhs_array_muxed;
						end
						9'd299: begin
							mem_ctrl_memorycontroller307 <= verilog_output_f_lhs_array_muxed;
						end
						9'd300: begin
							mem_ctrl_memorycontroller308 <= verilog_output_f_lhs_array_muxed;
						end
						9'd301: begin
							mem_ctrl_memorycontroller309 <= verilog_output_f_lhs_array_muxed;
						end
						9'd302: begin
							mem_ctrl_memorycontroller310 <= verilog_output_f_lhs_array_muxed;
						end
						9'd303: begin
							mem_ctrl_memorycontroller311 <= verilog_output_f_lhs_array_muxed;
						end
						9'd304: begin
							mem_ctrl_memorycontroller312 <= verilog_output_f_lhs_array_muxed;
						end
						9'd305: begin
							mem_ctrl_memorycontroller313 <= verilog_output_f_lhs_array_muxed;
						end
						9'd306: begin
							mem_ctrl_memorycontroller314 <= verilog_output_f_lhs_array_muxed;
						end
						9'd307: begin
							mem_ctrl_memorycontroller315 <= verilog_output_f_lhs_array_muxed;
						end
						9'd308: begin
							mem_ctrl_memorycontroller316 <= verilog_output_f_lhs_array_muxed;
						end
						9'd309: begin
							mem_ctrl_memorycontroller317 <= verilog_output_f_lhs_array_muxed;
						end
						9'd310: begin
							mem_ctrl_memorycontroller318 <= verilog_output_f_lhs_array_muxed;
						end
						9'd311: begin
							mem_ctrl_memorycontroller319 <= verilog_output_f_lhs_array_muxed;
						end
						9'd312: begin
							mem_ctrl_memorycontroller320 <= verilog_output_f_lhs_array_muxed;
						end
						9'd313: begin
							mem_ctrl_memorycontroller321 <= verilog_output_f_lhs_array_muxed;
						end
						9'd314: begin
							mem_ctrl_memorycontroller322 <= verilog_output_f_lhs_array_muxed;
						end
						9'd315: begin
							mem_ctrl_memorycontroller323 <= verilog_output_f_lhs_array_muxed;
						end
						9'd316: begin
							mem_ctrl_memorycontroller324 <= verilog_output_f_lhs_array_muxed;
						end
						9'd317: begin
							mem_ctrl_memorycontroller325 <= verilog_output_f_lhs_array_muxed;
						end
						9'd318: begin
							mem_ctrl_memorycontroller326 <= verilog_output_f_lhs_array_muxed;
						end
						9'd319: begin
							mem_ctrl_memorycontroller327 <= verilog_output_f_lhs_array_muxed;
						end
						9'd320: begin
							mem_ctrl_memorycontroller328 <= verilog_output_f_lhs_array_muxed;
						end
						9'd321: begin
							mem_ctrl_memorycontroller329 <= verilog_output_f_lhs_array_muxed;
						end
						9'd322: begin
							mem_ctrl_memorycontroller330 <= verilog_output_f_lhs_array_muxed;
						end
						9'd323: begin
							mem_ctrl_memorycontroller331 <= verilog_output_f_lhs_array_muxed;
						end
						9'd324: begin
							mem_ctrl_memorycontroller332 <= verilog_output_f_lhs_array_muxed;
						end
						9'd325: begin
							mem_ctrl_memorycontroller333 <= verilog_output_f_lhs_array_muxed;
						end
						9'd326: begin
							mem_ctrl_memorycontroller334 <= verilog_output_f_lhs_array_muxed;
						end
						9'd327: begin
							mem_ctrl_memorycontroller335 <= verilog_output_f_lhs_array_muxed;
						end
						9'd328: begin
							mem_ctrl_memorycontroller336 <= verilog_output_f_lhs_array_muxed;
						end
						9'd329: begin
							mem_ctrl_memorycontroller337 <= verilog_output_f_lhs_array_muxed;
						end
						9'd330: begin
							mem_ctrl_memorycontroller338 <= verilog_output_f_lhs_array_muxed;
						end
						9'd331: begin
							mem_ctrl_memorycontroller339 <= verilog_output_f_lhs_array_muxed;
						end
						9'd332: begin
							mem_ctrl_memorycontroller340 <= verilog_output_f_lhs_array_muxed;
						end
						9'd333: begin
							mem_ctrl_memorycontroller341 <= verilog_output_f_lhs_array_muxed;
						end
						9'd334: begin
							mem_ctrl_memorycontroller342 <= verilog_output_f_lhs_array_muxed;
						end
						9'd335: begin
							mem_ctrl_memorycontroller343 <= verilog_output_f_lhs_array_muxed;
						end
						9'd336: begin
							mem_ctrl_memorycontroller344 <= verilog_output_f_lhs_array_muxed;
						end
						9'd337: begin
							mem_ctrl_memorycontroller345 <= verilog_output_f_lhs_array_muxed;
						end
						9'd338: begin
							mem_ctrl_memorycontroller346 <= verilog_output_f_lhs_array_muxed;
						end
						9'd339: begin
							mem_ctrl_memorycontroller347 <= verilog_output_f_lhs_array_muxed;
						end
						9'd340: begin
							mem_ctrl_memorycontroller348 <= verilog_output_f_lhs_array_muxed;
						end
						9'd341: begin
							mem_ctrl_memorycontroller349 <= verilog_output_f_lhs_array_muxed;
						end
						9'd342: begin
							mem_ctrl_memorycontroller350 <= verilog_output_f_lhs_array_muxed;
						end
						9'd343: begin
							mem_ctrl_memorycontroller351 <= verilog_output_f_lhs_array_muxed;
						end
						9'd344: begin
							mem_ctrl_memorycontroller352 <= verilog_output_f_lhs_array_muxed;
						end
						9'd345: begin
							mem_ctrl_memorycontroller353 <= verilog_output_f_lhs_array_muxed;
						end
						9'd346: begin
							mem_ctrl_memorycontroller354 <= verilog_output_f_lhs_array_muxed;
						end
						9'd347: begin
							mem_ctrl_memorycontroller355 <= verilog_output_f_lhs_array_muxed;
						end
						9'd348: begin
							mem_ctrl_memorycontroller356 <= verilog_output_f_lhs_array_muxed;
						end
						9'd349: begin
							mem_ctrl_memorycontroller357 <= verilog_output_f_lhs_array_muxed;
						end
						9'd350: begin
							mem_ctrl_memorycontroller358 <= verilog_output_f_lhs_array_muxed;
						end
						9'd351: begin
							mem_ctrl_memorycontroller359 <= verilog_output_f_lhs_array_muxed;
						end
						9'd352: begin
							mem_ctrl_memorycontroller360 <= verilog_output_f_lhs_array_muxed;
						end
						9'd353: begin
							mem_ctrl_memorycontroller361 <= verilog_output_f_lhs_array_muxed;
						end
						9'd354: begin
							mem_ctrl_memorycontroller362 <= verilog_output_f_lhs_array_muxed;
						end
						9'd355: begin
							mem_ctrl_memorycontroller363 <= verilog_output_f_lhs_array_muxed;
						end
						9'd356: begin
							mem_ctrl_memorycontroller364 <= verilog_output_f_lhs_array_muxed;
						end
						9'd357: begin
							mem_ctrl_memorycontroller365 <= verilog_output_f_lhs_array_muxed;
						end
						9'd358: begin
							mem_ctrl_memorycontroller366 <= verilog_output_f_lhs_array_muxed;
						end
						9'd359: begin
							mem_ctrl_memorycontroller367 <= verilog_output_f_lhs_array_muxed;
						end
						9'd360: begin
							mem_ctrl_memorycontroller368 <= verilog_output_f_lhs_array_muxed;
						end
						9'd361: begin
							mem_ctrl_memorycontroller369 <= verilog_output_f_lhs_array_muxed;
						end
						9'd362: begin
							mem_ctrl_memorycontroller370 <= verilog_output_f_lhs_array_muxed;
						end
						9'd363: begin
							mem_ctrl_memorycontroller371 <= verilog_output_f_lhs_array_muxed;
						end
						9'd364: begin
							mem_ctrl_memorycontroller372 <= verilog_output_f_lhs_array_muxed;
						end
						9'd365: begin
							mem_ctrl_memorycontroller373 <= verilog_output_f_lhs_array_muxed;
						end
						9'd366: begin
							mem_ctrl_memorycontroller374 <= verilog_output_f_lhs_array_muxed;
						end
						9'd367: begin
							mem_ctrl_memorycontroller375 <= verilog_output_f_lhs_array_muxed;
						end
						9'd368: begin
							mem_ctrl_memorycontroller376 <= verilog_output_f_lhs_array_muxed;
						end
						9'd369: begin
							mem_ctrl_memorycontroller377 <= verilog_output_f_lhs_array_muxed;
						end
						9'd370: begin
							mem_ctrl_memorycontroller378 <= verilog_output_f_lhs_array_muxed;
						end
						9'd371: begin
							mem_ctrl_memorycontroller379 <= verilog_output_f_lhs_array_muxed;
						end
						9'd372: begin
							mem_ctrl_memorycontroller380 <= verilog_output_f_lhs_array_muxed;
						end
						9'd373: begin
							mem_ctrl_memorycontroller381 <= verilog_output_f_lhs_array_muxed;
						end
						9'd374: begin
							mem_ctrl_memorycontroller382 <= verilog_output_f_lhs_array_muxed;
						end
						9'd375: begin
							mem_ctrl_memorycontroller383 <= verilog_output_f_lhs_array_muxed;
						end
						9'd376: begin
							mem_ctrl_memorycontroller384 <= verilog_output_f_lhs_array_muxed;
						end
						9'd377: begin
							mem_ctrl_memorycontroller385 <= verilog_output_f_lhs_array_muxed;
						end
						9'd378: begin
							mem_ctrl_memorycontroller386 <= verilog_output_f_lhs_array_muxed;
						end
						9'd379: begin
							mem_ctrl_memorycontroller387 <= verilog_output_f_lhs_array_muxed;
						end
						9'd380: begin
							mem_ctrl_memorycontroller388 <= verilog_output_f_lhs_array_muxed;
						end
						9'd381: begin
							mem_ctrl_memorycontroller389 <= verilog_output_f_lhs_array_muxed;
						end
						9'd382: begin
							mem_ctrl_memorycontroller390 <= verilog_output_f_lhs_array_muxed;
						end
						9'd383: begin
							mem_ctrl_memorycontroller391 <= verilog_output_f_lhs_array_muxed;
						end
						9'd384: begin
							mem_ctrl_memorycontroller392 <= verilog_output_f_lhs_array_muxed;
						end
						9'd385: begin
							mem_ctrl_memorycontroller393 <= verilog_output_f_lhs_array_muxed;
						end
						9'd386: begin
							mem_ctrl_memorycontroller394 <= verilog_output_f_lhs_array_muxed;
						end
						9'd387: begin
							mem_ctrl_memorycontroller395 <= verilog_output_f_lhs_array_muxed;
						end
						9'd388: begin
							mem_ctrl_memorycontroller396 <= verilog_output_f_lhs_array_muxed;
						end
						9'd389: begin
							mem_ctrl_memorycontroller397 <= verilog_output_f_lhs_array_muxed;
						end
						9'd390: begin
							mem_ctrl_memorycontroller398 <= verilog_output_f_lhs_array_muxed;
						end
						9'd391: begin
							mem_ctrl_memorycontroller399 <= verilog_output_f_lhs_array_muxed;
						end
						9'd392: begin
							mem_ctrl_memorycontroller400 <= verilog_output_f_lhs_array_muxed;
						end
						9'd393: begin
							mem_ctrl_memorycontroller401 <= verilog_output_f_lhs_array_muxed;
						end
						9'd394: begin
							mem_ctrl_memorycontroller402 <= verilog_output_f_lhs_array_muxed;
						end
						9'd395: begin
							mem_ctrl_memorycontroller403 <= verilog_output_f_lhs_array_muxed;
						end
						9'd396: begin
							mem_ctrl_memorycontroller404 <= verilog_output_f_lhs_array_muxed;
						end
						9'd397: begin
							mem_ctrl_memorycontroller405 <= verilog_output_f_lhs_array_muxed;
						end
						9'd398: begin
							mem_ctrl_memorycontroller406 <= verilog_output_f_lhs_array_muxed;
						end
						9'd399: begin
							mem_ctrl_memorycontroller407 <= verilog_output_f_lhs_array_muxed;
						end
						9'd400: begin
							mem_ctrl_memorycontroller408 <= verilog_output_f_lhs_array_muxed;
						end
						9'd401: begin
							mem_ctrl_memorycontroller409 <= verilog_output_f_lhs_array_muxed;
						end
						9'd402: begin
							mem_ctrl_memorycontroller410 <= verilog_output_f_lhs_array_muxed;
						end
						9'd403: begin
							mem_ctrl_memorycontroller411 <= verilog_output_f_lhs_array_muxed;
						end
						9'd404: begin
							mem_ctrl_memorycontroller412 <= verilog_output_f_lhs_array_muxed;
						end
						9'd405: begin
							mem_ctrl_memorycontroller413 <= verilog_output_f_lhs_array_muxed;
						end
						9'd406: begin
							mem_ctrl_memorycontroller414 <= verilog_output_f_lhs_array_muxed;
						end
						9'd407: begin
							mem_ctrl_memorycontroller415 <= verilog_output_f_lhs_array_muxed;
						end
						9'd408: begin
							mem_ctrl_memorycontroller416 <= verilog_output_f_lhs_array_muxed;
						end
						9'd409: begin
							mem_ctrl_memorycontroller417 <= verilog_output_f_lhs_array_muxed;
						end
						9'd410: begin
							mem_ctrl_memorycontroller418 <= verilog_output_f_lhs_array_muxed;
						end
						9'd411: begin
							mem_ctrl_memorycontroller419 <= verilog_output_f_lhs_array_muxed;
						end
						9'd412: begin
							mem_ctrl_memorycontroller420 <= verilog_output_f_lhs_array_muxed;
						end
						9'd413: begin
							mem_ctrl_memorycontroller421 <= verilog_output_f_lhs_array_muxed;
						end
						9'd414: begin
							mem_ctrl_memorycontroller422 <= verilog_output_f_lhs_array_muxed;
						end
						9'd415: begin
							mem_ctrl_memorycontroller423 <= verilog_output_f_lhs_array_muxed;
						end
						9'd416: begin
							mem_ctrl_memorycontroller424 <= verilog_output_f_lhs_array_muxed;
						end
						9'd417: begin
							mem_ctrl_memorycontroller425 <= verilog_output_f_lhs_array_muxed;
						end
						9'd418: begin
							mem_ctrl_memorycontroller426 <= verilog_output_f_lhs_array_muxed;
						end
						9'd419: begin
							mem_ctrl_memorycontroller427 <= verilog_output_f_lhs_array_muxed;
						end
						9'd420: begin
							mem_ctrl_memorycontroller428 <= verilog_output_f_lhs_array_muxed;
						end
						9'd421: begin
							mem_ctrl_memorycontroller429 <= verilog_output_f_lhs_array_muxed;
						end
						9'd422: begin
							mem_ctrl_memorycontroller430 <= verilog_output_f_lhs_array_muxed;
						end
						9'd423: begin
							mem_ctrl_memorycontroller431 <= verilog_output_f_lhs_array_muxed;
						end
						9'd424: begin
							mem_ctrl_memorycontroller432 <= verilog_output_f_lhs_array_muxed;
						end
						9'd425: begin
							mem_ctrl_memorycontroller433 <= verilog_output_f_lhs_array_muxed;
						end
						9'd426: begin
							mem_ctrl_memorycontroller434 <= verilog_output_f_lhs_array_muxed;
						end
						9'd427: begin
							mem_ctrl_memorycontroller435 <= verilog_output_f_lhs_array_muxed;
						end
						9'd428: begin
							mem_ctrl_memorycontroller436 <= verilog_output_f_lhs_array_muxed;
						end
						9'd429: begin
							mem_ctrl_memorycontroller437 <= verilog_output_f_lhs_array_muxed;
						end
						9'd430: begin
							mem_ctrl_memorycontroller438 <= verilog_output_f_lhs_array_muxed;
						end
						9'd431: begin
							mem_ctrl_memorycontroller439 <= verilog_output_f_lhs_array_muxed;
						end
						9'd432: begin
							mem_ctrl_memorycontroller440 <= verilog_output_f_lhs_array_muxed;
						end
						9'd433: begin
							mem_ctrl_memorycontroller441 <= verilog_output_f_lhs_array_muxed;
						end
						9'd434: begin
							mem_ctrl_memorycontroller442 <= verilog_output_f_lhs_array_muxed;
						end
						9'd435: begin
							mem_ctrl_memorycontroller443 <= verilog_output_f_lhs_array_muxed;
						end
						9'd436: begin
							mem_ctrl_memorycontroller444 <= verilog_output_f_lhs_array_muxed;
						end
						9'd437: begin
							mem_ctrl_memorycontroller445 <= verilog_output_f_lhs_array_muxed;
						end
						9'd438: begin
							mem_ctrl_memorycontroller446 <= verilog_output_f_lhs_array_muxed;
						end
						9'd439: begin
							mem_ctrl_memorycontroller447 <= verilog_output_f_lhs_array_muxed;
						end
						9'd440: begin
							mem_ctrl_memorycontroller448 <= verilog_output_f_lhs_array_muxed;
						end
						9'd441: begin
							mem_ctrl_memorycontroller449 <= verilog_output_f_lhs_array_muxed;
						end
						9'd442: begin
							mem_ctrl_memorycontroller450 <= verilog_output_f_lhs_array_muxed;
						end
						9'd443: begin
							mem_ctrl_memorycontroller451 <= verilog_output_f_lhs_array_muxed;
						end
						9'd444: begin
							mem_ctrl_memorycontroller452 <= verilog_output_f_lhs_array_muxed;
						end
						9'd445: begin
							mem_ctrl_memorycontroller453 <= verilog_output_f_lhs_array_muxed;
						end
						9'd446: begin
							mem_ctrl_memorycontroller454 <= verilog_output_f_lhs_array_muxed;
						end
						9'd447: begin
							mem_ctrl_memorycontroller455 <= verilog_output_f_lhs_array_muxed;
						end
						9'd448: begin
							mem_ctrl_memorycontroller456 <= verilog_output_f_lhs_array_muxed;
						end
						9'd449: begin
							mem_ctrl_memorycontroller457 <= verilog_output_f_lhs_array_muxed;
						end
						9'd450: begin
							mem_ctrl_memorycontroller458 <= verilog_output_f_lhs_array_muxed;
						end
						9'd451: begin
							mem_ctrl_memorycontroller459 <= verilog_output_f_lhs_array_muxed;
						end
						9'd452: begin
							mem_ctrl_memorycontroller460 <= verilog_output_f_lhs_array_muxed;
						end
						9'd453: begin
							mem_ctrl_memorycontroller461 <= verilog_output_f_lhs_array_muxed;
						end
						9'd454: begin
							mem_ctrl_memorycontroller462 <= verilog_output_f_lhs_array_muxed;
						end
						9'd455: begin
							mem_ctrl_memorycontroller463 <= verilog_output_f_lhs_array_muxed;
						end
						9'd456: begin
							mem_ctrl_memorycontroller464 <= verilog_output_f_lhs_array_muxed;
						end
						9'd457: begin
							mem_ctrl_memorycontroller465 <= verilog_output_f_lhs_array_muxed;
						end
						9'd458: begin
							mem_ctrl_memorycontroller466 <= verilog_output_f_lhs_array_muxed;
						end
						9'd459: begin
							mem_ctrl_memorycontroller467 <= verilog_output_f_lhs_array_muxed;
						end
						9'd460: begin
							mem_ctrl_memorycontroller468 <= verilog_output_f_lhs_array_muxed;
						end
						9'd461: begin
							mem_ctrl_memorycontroller469 <= verilog_output_f_lhs_array_muxed;
						end
						9'd462: begin
							mem_ctrl_memorycontroller470 <= verilog_output_f_lhs_array_muxed;
						end
						9'd463: begin
							mem_ctrl_memorycontroller471 <= verilog_output_f_lhs_array_muxed;
						end
						9'd464: begin
							mem_ctrl_memorycontroller472 <= verilog_output_f_lhs_array_muxed;
						end
						9'd465: begin
							mem_ctrl_memorycontroller473 <= verilog_output_f_lhs_array_muxed;
						end
						9'd466: begin
							mem_ctrl_memorycontroller474 <= verilog_output_f_lhs_array_muxed;
						end
						9'd467: begin
							mem_ctrl_memorycontroller475 <= verilog_output_f_lhs_array_muxed;
						end
						9'd468: begin
							mem_ctrl_memorycontroller476 <= verilog_output_f_lhs_array_muxed;
						end
						9'd469: begin
							mem_ctrl_memorycontroller477 <= verilog_output_f_lhs_array_muxed;
						end
						9'd470: begin
							mem_ctrl_memorycontroller478 <= verilog_output_f_lhs_array_muxed;
						end
						9'd471: begin
							mem_ctrl_memorycontroller479 <= verilog_output_f_lhs_array_muxed;
						end
						9'd472: begin
							mem_ctrl_memorycontroller480 <= verilog_output_f_lhs_array_muxed;
						end
						9'd473: begin
							mem_ctrl_memorycontroller481 <= verilog_output_f_lhs_array_muxed;
						end
						9'd474: begin
							mem_ctrl_memorycontroller482 <= verilog_output_f_lhs_array_muxed;
						end
						9'd475: begin
							mem_ctrl_memorycontroller483 <= verilog_output_f_lhs_array_muxed;
						end
						9'd476: begin
							mem_ctrl_memorycontroller484 <= verilog_output_f_lhs_array_muxed;
						end
						9'd477: begin
							mem_ctrl_memorycontroller485 <= verilog_output_f_lhs_array_muxed;
						end
						9'd478: begin
							mem_ctrl_memorycontroller486 <= verilog_output_f_lhs_array_muxed;
						end
						9'd479: begin
							mem_ctrl_memorycontroller487 <= verilog_output_f_lhs_array_muxed;
						end
						9'd480: begin
							mem_ctrl_memorycontroller488 <= verilog_output_f_lhs_array_muxed;
						end
						9'd481: begin
							mem_ctrl_memorycontroller489 <= verilog_output_f_lhs_array_muxed;
						end
						9'd482: begin
							mem_ctrl_memorycontroller490 <= verilog_output_f_lhs_array_muxed;
						end
						9'd483: begin
							mem_ctrl_memorycontroller491 <= verilog_output_f_lhs_array_muxed;
						end
						9'd484: begin
							mem_ctrl_memorycontroller492 <= verilog_output_f_lhs_array_muxed;
						end
						9'd485: begin
							mem_ctrl_memorycontroller493 <= verilog_output_f_lhs_array_muxed;
						end
						9'd486: begin
							mem_ctrl_memorycontroller494 <= verilog_output_f_lhs_array_muxed;
						end
						9'd487: begin
							mem_ctrl_memorycontroller495 <= verilog_output_f_lhs_array_muxed;
						end
						9'd488: begin
							mem_ctrl_memorycontroller496 <= verilog_output_f_lhs_array_muxed;
						end
						9'd489: begin
							mem_ctrl_memorycontroller497 <= verilog_output_f_lhs_array_muxed;
						end
						9'd490: begin
							mem_ctrl_memorycontroller498 <= verilog_output_f_lhs_array_muxed;
						end
						9'd491: begin
							mem_ctrl_memorycontroller499 <= verilog_output_f_lhs_array_muxed;
						end
						9'd492: begin
							mem_ctrl_memorycontroller500 <= verilog_output_f_lhs_array_muxed;
						end
						9'd493: begin
							mem_ctrl_memorycontroller501 <= verilog_output_f_lhs_array_muxed;
						end
						9'd494: begin
							mem_ctrl_memorycontroller502 <= verilog_output_f_lhs_array_muxed;
						end
						9'd495: begin
							mem_ctrl_memorycontroller503 <= verilog_output_f_lhs_array_muxed;
						end
						9'd496: begin
							mem_ctrl_memorycontroller504 <= verilog_output_f_lhs_array_muxed;
						end
						9'd497: begin
							mem_ctrl_memorycontroller505 <= verilog_output_f_lhs_array_muxed;
						end
						9'd498: begin
							mem_ctrl_memorycontroller506 <= verilog_output_f_lhs_array_muxed;
						end
						9'd499: begin
							mem_ctrl_memorycontroller507 <= verilog_output_f_lhs_array_muxed;
						end
						9'd500: begin
							mem_ctrl_memorycontroller508 <= verilog_output_f_lhs_array_muxed;
						end
						9'd501: begin
							mem_ctrl_memorycontroller509 <= verilog_output_f_lhs_array_muxed;
						end
						9'd502: begin
							mem_ctrl_memorycontroller510 <= verilog_output_f_lhs_array_muxed;
						end
						9'd503: begin
							mem_ctrl_memorycontroller511 <= verilog_output_f_lhs_array_muxed;
						end
						9'd504: begin
							mem_ctrl_memorycontroller512 <= verilog_output_f_lhs_array_muxed;
						end
						9'd505: begin
							mem_ctrl_memorycontroller513 <= verilog_output_f_lhs_array_muxed;
						end
						9'd506: begin
							mem_ctrl_memorycontroller514 <= verilog_output_f_lhs_array_muxed;
						end
						9'd507: begin
							mem_ctrl_memorycontroller515 <= verilog_output_f_lhs_array_muxed;
						end
						9'd508: begin
							mem_ctrl_memorycontroller516 <= verilog_output_f_lhs_array_muxed;
						end
						9'd509: begin
							mem_ctrl_memorycontroller517 <= verilog_output_f_lhs_array_muxed;
						end
						9'd510: begin
							mem_ctrl_memorycontroller518 <= verilog_output_f_lhs_array_muxed;
						end
						9'd511: begin
							mem_ctrl_memorycontroller519 <= verilog_output_f_lhs_array_muxed;
						end
						10'd512: begin
							mem_ctrl_memorycontroller520 <= verilog_output_f_lhs_array_muxed;
						end
						10'd513: begin
							mem_ctrl_memorycontroller521 <= verilog_output_f_lhs_array_muxed;
						end
						10'd514: begin
							mem_ctrl_memorycontroller522 <= verilog_output_f_lhs_array_muxed;
						end
						10'd515: begin
							mem_ctrl_memorycontroller523 <= verilog_output_f_lhs_array_muxed;
						end
						10'd516: begin
							mem_ctrl_memorycontroller524 <= verilog_output_f_lhs_array_muxed;
						end
						10'd517: begin
							mem_ctrl_memorycontroller525 <= verilog_output_f_lhs_array_muxed;
						end
						10'd518: begin
							mem_ctrl_memorycontroller526 <= verilog_output_f_lhs_array_muxed;
						end
						10'd519: begin
							mem_ctrl_memorycontroller527 <= verilog_output_f_lhs_array_muxed;
						end
						10'd520: begin
							mem_ctrl_memorycontroller528 <= verilog_output_f_lhs_array_muxed;
						end
						10'd521: begin
							mem_ctrl_memorycontroller529 <= verilog_output_f_lhs_array_muxed;
						end
						10'd522: begin
							mem_ctrl_memorycontroller530 <= verilog_output_f_lhs_array_muxed;
						end
						10'd523: begin
							mem_ctrl_memorycontroller531 <= verilog_output_f_lhs_array_muxed;
						end
						10'd524: begin
							mem_ctrl_memorycontroller532 <= verilog_output_f_lhs_array_muxed;
						end
						10'd525: begin
							mem_ctrl_memorycontroller533 <= verilog_output_f_lhs_array_muxed;
						end
						10'd526: begin
							mem_ctrl_memorycontroller534 <= verilog_output_f_lhs_array_muxed;
						end
						10'd527: begin
							mem_ctrl_memorycontroller535 <= verilog_output_f_lhs_array_muxed;
						end
						10'd528: begin
							mem_ctrl_memorycontroller536 <= verilog_output_f_lhs_array_muxed;
						end
						10'd529: begin
							mem_ctrl_memorycontroller537 <= verilog_output_f_lhs_array_muxed;
						end
						10'd530: begin
							mem_ctrl_memorycontroller538 <= verilog_output_f_lhs_array_muxed;
						end
						10'd531: begin
							mem_ctrl_memorycontroller539 <= verilog_output_f_lhs_array_muxed;
						end
						10'd532: begin
							mem_ctrl_memorycontroller540 <= verilog_output_f_lhs_array_muxed;
						end
						10'd533: begin
							mem_ctrl_memorycontroller541 <= verilog_output_f_lhs_array_muxed;
						end
						10'd534: begin
							mem_ctrl_memorycontroller542 <= verilog_output_f_lhs_array_muxed;
						end
						10'd535: begin
							mem_ctrl_memorycontroller543 <= verilog_output_f_lhs_array_muxed;
						end
						10'd536: begin
							mem_ctrl_memorycontroller544 <= verilog_output_f_lhs_array_muxed;
						end
						10'd537: begin
							mem_ctrl_memorycontroller545 <= verilog_output_f_lhs_array_muxed;
						end
						10'd538: begin
							mem_ctrl_memorycontroller546 <= verilog_output_f_lhs_array_muxed;
						end
						10'd539: begin
							mem_ctrl_memorycontroller547 <= verilog_output_f_lhs_array_muxed;
						end
						10'd540: begin
							mem_ctrl_memorycontroller548 <= verilog_output_f_lhs_array_muxed;
						end
						10'd541: begin
							mem_ctrl_memorycontroller549 <= verilog_output_f_lhs_array_muxed;
						end
						10'd542: begin
							mem_ctrl_memorycontroller550 <= verilog_output_f_lhs_array_muxed;
						end
						10'd543: begin
							mem_ctrl_memorycontroller551 <= verilog_output_f_lhs_array_muxed;
						end
						10'd544: begin
							mem_ctrl_memorycontroller552 <= verilog_output_f_lhs_array_muxed;
						end
						10'd545: begin
							mem_ctrl_memorycontroller553 <= verilog_output_f_lhs_array_muxed;
						end
						10'd546: begin
							mem_ctrl_memorycontroller554 <= verilog_output_f_lhs_array_muxed;
						end
						10'd547: begin
							mem_ctrl_memorycontroller555 <= verilog_output_f_lhs_array_muxed;
						end
						10'd548: begin
							mem_ctrl_memorycontroller556 <= verilog_output_f_lhs_array_muxed;
						end
						10'd549: begin
							mem_ctrl_memorycontroller557 <= verilog_output_f_lhs_array_muxed;
						end
						10'd550: begin
							mem_ctrl_memorycontroller558 <= verilog_output_f_lhs_array_muxed;
						end
						10'd551: begin
							mem_ctrl_memorycontroller559 <= verilog_output_f_lhs_array_muxed;
						end
						10'd552: begin
							mem_ctrl_memorycontroller560 <= verilog_output_f_lhs_array_muxed;
						end
						10'd553: begin
							mem_ctrl_memorycontroller561 <= verilog_output_f_lhs_array_muxed;
						end
						10'd554: begin
							mem_ctrl_memorycontroller562 <= verilog_output_f_lhs_array_muxed;
						end
						10'd555: begin
							mem_ctrl_memorycontroller563 <= verilog_output_f_lhs_array_muxed;
						end
						10'd556: begin
							mem_ctrl_memorycontroller564 <= verilog_output_f_lhs_array_muxed;
						end
						10'd557: begin
							mem_ctrl_memorycontroller565 <= verilog_output_f_lhs_array_muxed;
						end
						10'd558: begin
							mem_ctrl_memorycontroller566 <= verilog_output_f_lhs_array_muxed;
						end
						10'd559: begin
							mem_ctrl_memorycontroller567 <= verilog_output_f_lhs_array_muxed;
						end
						10'd560: begin
							mem_ctrl_memorycontroller568 <= verilog_output_f_lhs_array_muxed;
						end
						10'd561: begin
							mem_ctrl_memorycontroller569 <= verilog_output_f_lhs_array_muxed;
						end
						10'd562: begin
							mem_ctrl_memorycontroller570 <= verilog_output_f_lhs_array_muxed;
						end
						10'd563: begin
							mem_ctrl_memorycontroller571 <= verilog_output_f_lhs_array_muxed;
						end
						10'd564: begin
							mem_ctrl_memorycontroller572 <= verilog_output_f_lhs_array_muxed;
						end
						10'd565: begin
							mem_ctrl_memorycontroller573 <= verilog_output_f_lhs_array_muxed;
						end
						10'd566: begin
							mem_ctrl_memorycontroller574 <= verilog_output_f_lhs_array_muxed;
						end
						10'd567: begin
							mem_ctrl_memorycontroller575 <= verilog_output_f_lhs_array_muxed;
						end
						10'd568: begin
							mem_ctrl_memorycontroller576 <= verilog_output_f_lhs_array_muxed;
						end
						10'd569: begin
							mem_ctrl_memorycontroller577 <= verilog_output_f_lhs_array_muxed;
						end
						10'd570: begin
							mem_ctrl_memorycontroller578 <= verilog_output_f_lhs_array_muxed;
						end
						10'd571: begin
							mem_ctrl_memorycontroller579 <= verilog_output_f_lhs_array_muxed;
						end
						10'd572: begin
							mem_ctrl_memorycontroller580 <= verilog_output_f_lhs_array_muxed;
						end
						10'd573: begin
							mem_ctrl_memorycontroller581 <= verilog_output_f_lhs_array_muxed;
						end
						10'd574: begin
							mem_ctrl_memorycontroller582 <= verilog_output_f_lhs_array_muxed;
						end
						10'd575: begin
							mem_ctrl_memorycontroller583 <= verilog_output_f_lhs_array_muxed;
						end
						10'd576: begin
							mem_ctrl_memorycontroller584 <= verilog_output_f_lhs_array_muxed;
						end
						10'd577: begin
							mem_ctrl_memorycontroller585 <= verilog_output_f_lhs_array_muxed;
						end
						10'd578: begin
							mem_ctrl_memorycontroller586 <= verilog_output_f_lhs_array_muxed;
						end
						10'd579: begin
							mem_ctrl_memorycontroller587 <= verilog_output_f_lhs_array_muxed;
						end
						10'd580: begin
							mem_ctrl_memorycontroller588 <= verilog_output_f_lhs_array_muxed;
						end
						10'd581: begin
							mem_ctrl_memorycontroller589 <= verilog_output_f_lhs_array_muxed;
						end
						10'd582: begin
							mem_ctrl_memorycontroller590 <= verilog_output_f_lhs_array_muxed;
						end
						10'd583: begin
							mem_ctrl_memorycontroller591 <= verilog_output_f_lhs_array_muxed;
						end
						10'd584: begin
							mem_ctrl_memorycontroller592 <= verilog_output_f_lhs_array_muxed;
						end
						10'd585: begin
							mem_ctrl_memorycontroller593 <= verilog_output_f_lhs_array_muxed;
						end
						10'd586: begin
							mem_ctrl_memorycontroller594 <= verilog_output_f_lhs_array_muxed;
						end
						10'd587: begin
							mem_ctrl_memorycontroller595 <= verilog_output_f_lhs_array_muxed;
						end
						10'd588: begin
							mem_ctrl_memorycontroller596 <= verilog_output_f_lhs_array_muxed;
						end
						10'd589: begin
							mem_ctrl_memorycontroller597 <= verilog_output_f_lhs_array_muxed;
						end
						10'd590: begin
							mem_ctrl_memorycontroller598 <= verilog_output_f_lhs_array_muxed;
						end
						10'd591: begin
							mem_ctrl_memorycontroller599 <= verilog_output_f_lhs_array_muxed;
						end
						10'd592: begin
							mem_ctrl_memorycontroller600 <= verilog_output_f_lhs_array_muxed;
						end
						10'd593: begin
							mem_ctrl_memorycontroller601 <= verilog_output_f_lhs_array_muxed;
						end
						10'd594: begin
							mem_ctrl_memorycontroller602 <= verilog_output_f_lhs_array_muxed;
						end
						10'd595: begin
							mem_ctrl_memorycontroller603 <= verilog_output_f_lhs_array_muxed;
						end
						10'd596: begin
							mem_ctrl_memorycontroller604 <= verilog_output_f_lhs_array_muxed;
						end
						10'd597: begin
							mem_ctrl_memorycontroller605 <= verilog_output_f_lhs_array_muxed;
						end
						10'd598: begin
							mem_ctrl_memorycontroller606 <= verilog_output_f_lhs_array_muxed;
						end
						10'd599: begin
							mem_ctrl_memorycontroller607 <= verilog_output_f_lhs_array_muxed;
						end
						10'd600: begin
							mem_ctrl_memorycontroller608 <= verilog_output_f_lhs_array_muxed;
						end
						10'd601: begin
							mem_ctrl_memorycontroller609 <= verilog_output_f_lhs_array_muxed;
						end
						10'd602: begin
							mem_ctrl_memorycontroller610 <= verilog_output_f_lhs_array_muxed;
						end
						10'd603: begin
							mem_ctrl_memorycontroller611 <= verilog_output_f_lhs_array_muxed;
						end
						10'd604: begin
							mem_ctrl_memorycontroller612 <= verilog_output_f_lhs_array_muxed;
						end
						10'd605: begin
							mem_ctrl_memorycontroller613 <= verilog_output_f_lhs_array_muxed;
						end
						10'd606: begin
							mem_ctrl_memorycontroller614 <= verilog_output_f_lhs_array_muxed;
						end
						10'd607: begin
							mem_ctrl_memorycontroller615 <= verilog_output_f_lhs_array_muxed;
						end
						10'd608: begin
							mem_ctrl_memorycontroller616 <= verilog_output_f_lhs_array_muxed;
						end
						10'd609: begin
							mem_ctrl_memorycontroller617 <= verilog_output_f_lhs_array_muxed;
						end
						10'd610: begin
							mem_ctrl_memorycontroller618 <= verilog_output_f_lhs_array_muxed;
						end
						10'd611: begin
							mem_ctrl_memorycontroller619 <= verilog_output_f_lhs_array_muxed;
						end
						10'd612: begin
							mem_ctrl_memorycontroller620 <= verilog_output_f_lhs_array_muxed;
						end
						10'd613: begin
							mem_ctrl_memorycontroller621 <= verilog_output_f_lhs_array_muxed;
						end
						10'd614: begin
							mem_ctrl_memorycontroller622 <= verilog_output_f_lhs_array_muxed;
						end
						10'd615: begin
							mem_ctrl_memorycontroller623 <= verilog_output_f_lhs_array_muxed;
						end
						10'd616: begin
							mem_ctrl_memorycontroller624 <= verilog_output_f_lhs_array_muxed;
						end
						10'd617: begin
							mem_ctrl_memorycontroller625 <= verilog_output_f_lhs_array_muxed;
						end
						10'd618: begin
							mem_ctrl_memorycontroller626 <= verilog_output_f_lhs_array_muxed;
						end
						10'd619: begin
							mem_ctrl_memorycontroller627 <= verilog_output_f_lhs_array_muxed;
						end
						10'd620: begin
							mem_ctrl_memorycontroller628 <= verilog_output_f_lhs_array_muxed;
						end
						10'd621: begin
							mem_ctrl_memorycontroller629 <= verilog_output_f_lhs_array_muxed;
						end
						10'd622: begin
							mem_ctrl_memorycontroller630 <= verilog_output_f_lhs_array_muxed;
						end
						10'd623: begin
							mem_ctrl_memorycontroller631 <= verilog_output_f_lhs_array_muxed;
						end
						10'd624: begin
							mem_ctrl_memorycontroller632 <= verilog_output_f_lhs_array_muxed;
						end
						10'd625: begin
							mem_ctrl_memorycontroller633 <= verilog_output_f_lhs_array_muxed;
						end
						10'd626: begin
							mem_ctrl_memorycontroller634 <= verilog_output_f_lhs_array_muxed;
						end
						10'd627: begin
							mem_ctrl_memorycontroller635 <= verilog_output_f_lhs_array_muxed;
						end
						10'd628: begin
							mem_ctrl_memorycontroller636 <= verilog_output_f_lhs_array_muxed;
						end
						10'd629: begin
							mem_ctrl_memorycontroller637 <= verilog_output_f_lhs_array_muxed;
						end
						10'd630: begin
							mem_ctrl_memorycontroller638 <= verilog_output_f_lhs_array_muxed;
						end
						10'd631: begin
							mem_ctrl_memorycontroller639 <= verilog_output_f_lhs_array_muxed;
						end
						10'd632: begin
							mem_ctrl_memorycontroller640 <= verilog_output_f_lhs_array_muxed;
						end
						10'd633: begin
							mem_ctrl_memorycontroller641 <= verilog_output_f_lhs_array_muxed;
						end
						10'd634: begin
							mem_ctrl_memorycontroller642 <= verilog_output_f_lhs_array_muxed;
						end
						10'd635: begin
							mem_ctrl_memorycontroller643 <= verilog_output_f_lhs_array_muxed;
						end
						10'd636: begin
							mem_ctrl_memorycontroller644 <= verilog_output_f_lhs_array_muxed;
						end
						10'd637: begin
							mem_ctrl_memorycontroller645 <= verilog_output_f_lhs_array_muxed;
						end
						10'd638: begin
							mem_ctrl_memorycontroller646 <= verilog_output_f_lhs_array_muxed;
						end
						10'd639: begin
							mem_ctrl_memorycontroller647 <= verilog_output_f_lhs_array_muxed;
						end
						10'd640: begin
							mem_ctrl_memorycontroller648 <= verilog_output_f_lhs_array_muxed;
						end
						10'd641: begin
							mem_ctrl_memorycontroller649 <= verilog_output_f_lhs_array_muxed;
						end
						10'd642: begin
							mem_ctrl_memorycontroller650 <= verilog_output_f_lhs_array_muxed;
						end
						10'd643: begin
							mem_ctrl_memorycontroller651 <= verilog_output_f_lhs_array_muxed;
						end
						10'd644: begin
							mem_ctrl_memorycontroller652 <= verilog_output_f_lhs_array_muxed;
						end
						10'd645: begin
							mem_ctrl_memorycontroller653 <= verilog_output_f_lhs_array_muxed;
						end
						10'd646: begin
							mem_ctrl_memorycontroller654 <= verilog_output_f_lhs_array_muxed;
						end
						10'd647: begin
							mem_ctrl_memorycontroller655 <= verilog_output_f_lhs_array_muxed;
						end
						10'd648: begin
							mem_ctrl_memorycontroller656 <= verilog_output_f_lhs_array_muxed;
						end
						10'd649: begin
							mem_ctrl_memorycontroller657 <= verilog_output_f_lhs_array_muxed;
						end
						10'd650: begin
							mem_ctrl_memorycontroller658 <= verilog_output_f_lhs_array_muxed;
						end
						10'd651: begin
							mem_ctrl_memorycontroller659 <= verilog_output_f_lhs_array_muxed;
						end
						10'd652: begin
							mem_ctrl_memorycontroller660 <= verilog_output_f_lhs_array_muxed;
						end
						10'd653: begin
							mem_ctrl_memorycontroller661 <= verilog_output_f_lhs_array_muxed;
						end
						10'd654: begin
							mem_ctrl_memorycontroller662 <= verilog_output_f_lhs_array_muxed;
						end
						10'd655: begin
							mem_ctrl_memorycontroller663 <= verilog_output_f_lhs_array_muxed;
						end
						10'd656: begin
							mem_ctrl_memorycontroller664 <= verilog_output_f_lhs_array_muxed;
						end
						10'd657: begin
							mem_ctrl_memorycontroller665 <= verilog_output_f_lhs_array_muxed;
						end
						10'd658: begin
							mem_ctrl_memorycontroller666 <= verilog_output_f_lhs_array_muxed;
						end
						10'd659: begin
							mem_ctrl_memorycontroller667 <= verilog_output_f_lhs_array_muxed;
						end
						10'd660: begin
							mem_ctrl_memorycontroller668 <= verilog_output_f_lhs_array_muxed;
						end
						10'd661: begin
							mem_ctrl_memorycontroller669 <= verilog_output_f_lhs_array_muxed;
						end
						10'd662: begin
							mem_ctrl_memorycontroller670 <= verilog_output_f_lhs_array_muxed;
						end
						10'd663: begin
							mem_ctrl_memorycontroller671 <= verilog_output_f_lhs_array_muxed;
						end
						10'd664: begin
							mem_ctrl_memorycontroller672 <= verilog_output_f_lhs_array_muxed;
						end
						10'd665: begin
							mem_ctrl_memorycontroller673 <= verilog_output_f_lhs_array_muxed;
						end
						10'd666: begin
							mem_ctrl_memorycontroller674 <= verilog_output_f_lhs_array_muxed;
						end
						10'd667: begin
							mem_ctrl_memorycontroller675 <= verilog_output_f_lhs_array_muxed;
						end
						10'd668: begin
							mem_ctrl_memorycontroller676 <= verilog_output_f_lhs_array_muxed;
						end
						10'd669: begin
							mem_ctrl_memorycontroller677 <= verilog_output_f_lhs_array_muxed;
						end
						10'd670: begin
							mem_ctrl_memorycontroller678 <= verilog_output_f_lhs_array_muxed;
						end
						10'd671: begin
							mem_ctrl_memorycontroller679 <= verilog_output_f_lhs_array_muxed;
						end
						10'd672: begin
							mem_ctrl_memorycontroller680 <= verilog_output_f_lhs_array_muxed;
						end
						10'd673: begin
							mem_ctrl_memorycontroller681 <= verilog_output_f_lhs_array_muxed;
						end
						10'd674: begin
							mem_ctrl_memorycontroller682 <= verilog_output_f_lhs_array_muxed;
						end
						10'd675: begin
							mem_ctrl_memorycontroller683 <= verilog_output_f_lhs_array_muxed;
						end
						10'd676: begin
							mem_ctrl_memorycontroller684 <= verilog_output_f_lhs_array_muxed;
						end
						10'd677: begin
							mem_ctrl_memorycontroller685 <= verilog_output_f_lhs_array_muxed;
						end
						10'd678: begin
							mem_ctrl_memorycontroller686 <= verilog_output_f_lhs_array_muxed;
						end
						10'd679: begin
							mem_ctrl_memorycontroller687 <= verilog_output_f_lhs_array_muxed;
						end
						10'd680: begin
							mem_ctrl_memorycontroller688 <= verilog_output_f_lhs_array_muxed;
						end
						10'd681: begin
							mem_ctrl_memorycontroller689 <= verilog_output_f_lhs_array_muxed;
						end
						10'd682: begin
							mem_ctrl_memorycontroller690 <= verilog_output_f_lhs_array_muxed;
						end
						10'd683: begin
							mem_ctrl_memorycontroller691 <= verilog_output_f_lhs_array_muxed;
						end
						10'd684: begin
							mem_ctrl_memorycontroller692 <= verilog_output_f_lhs_array_muxed;
						end
						10'd685: begin
							mem_ctrl_memorycontroller693 <= verilog_output_f_lhs_array_muxed;
						end
						10'd686: begin
							mem_ctrl_memorycontroller694 <= verilog_output_f_lhs_array_muxed;
						end
						10'd687: begin
							mem_ctrl_memorycontroller695 <= verilog_output_f_lhs_array_muxed;
						end
						10'd688: begin
							mem_ctrl_memorycontroller696 <= verilog_output_f_lhs_array_muxed;
						end
						10'd689: begin
							mem_ctrl_memorycontroller697 <= verilog_output_f_lhs_array_muxed;
						end
						10'd690: begin
							mem_ctrl_memorycontroller698 <= verilog_output_f_lhs_array_muxed;
						end
						10'd691: begin
							mem_ctrl_memorycontroller699 <= verilog_output_f_lhs_array_muxed;
						end
						10'd692: begin
							mem_ctrl_memorycontroller700 <= verilog_output_f_lhs_array_muxed;
						end
						10'd693: begin
							mem_ctrl_memorycontroller701 <= verilog_output_f_lhs_array_muxed;
						end
						10'd694: begin
							mem_ctrl_memorycontroller702 <= verilog_output_f_lhs_array_muxed;
						end
						10'd695: begin
							mem_ctrl_memorycontroller703 <= verilog_output_f_lhs_array_muxed;
						end
						10'd696: begin
							mem_ctrl_memorycontroller704 <= verilog_output_f_lhs_array_muxed;
						end
						10'd697: begin
							mem_ctrl_memorycontroller705 <= verilog_output_f_lhs_array_muxed;
						end
						10'd698: begin
							mem_ctrl_memorycontroller706 <= verilog_output_f_lhs_array_muxed;
						end
						10'd699: begin
							mem_ctrl_memorycontroller707 <= verilog_output_f_lhs_array_muxed;
						end
						10'd700: begin
							mem_ctrl_memorycontroller708 <= verilog_output_f_lhs_array_muxed;
						end
						10'd701: begin
							mem_ctrl_memorycontroller709 <= verilog_output_f_lhs_array_muxed;
						end
						10'd702: begin
							mem_ctrl_memorycontroller710 <= verilog_output_f_lhs_array_muxed;
						end
						10'd703: begin
							mem_ctrl_memorycontroller711 <= verilog_output_f_lhs_array_muxed;
						end
						10'd704: begin
							mem_ctrl_memorycontroller712 <= verilog_output_f_lhs_array_muxed;
						end
						10'd705: begin
							mem_ctrl_memorycontroller713 <= verilog_output_f_lhs_array_muxed;
						end
						10'd706: begin
							mem_ctrl_memorycontroller714 <= verilog_output_f_lhs_array_muxed;
						end
						10'd707: begin
							mem_ctrl_memorycontroller715 <= verilog_output_f_lhs_array_muxed;
						end
						10'd708: begin
							mem_ctrl_memorycontroller716 <= verilog_output_f_lhs_array_muxed;
						end
						10'd709: begin
							mem_ctrl_memorycontroller717 <= verilog_output_f_lhs_array_muxed;
						end
						10'd710: begin
							mem_ctrl_memorycontroller718 <= verilog_output_f_lhs_array_muxed;
						end
						10'd711: begin
							mem_ctrl_memorycontroller719 <= verilog_output_f_lhs_array_muxed;
						end
						10'd712: begin
							mem_ctrl_memorycontroller720 <= verilog_output_f_lhs_array_muxed;
						end
						10'd713: begin
							mem_ctrl_memorycontroller721 <= verilog_output_f_lhs_array_muxed;
						end
						10'd714: begin
							mem_ctrl_memorycontroller722 <= verilog_output_f_lhs_array_muxed;
						end
						10'd715: begin
							mem_ctrl_memorycontroller723 <= verilog_output_f_lhs_array_muxed;
						end
						10'd716: begin
							mem_ctrl_memorycontroller724 <= verilog_output_f_lhs_array_muxed;
						end
						10'd717: begin
							mem_ctrl_memorycontroller725 <= verilog_output_f_lhs_array_muxed;
						end
						10'd718: begin
							mem_ctrl_memorycontroller726 <= verilog_output_f_lhs_array_muxed;
						end
						10'd719: begin
							mem_ctrl_memorycontroller727 <= verilog_output_f_lhs_array_muxed;
						end
						10'd720: begin
							mem_ctrl_memorycontroller728 <= verilog_output_f_lhs_array_muxed;
						end
						10'd721: begin
							mem_ctrl_memorycontroller729 <= verilog_output_f_lhs_array_muxed;
						end
						10'd722: begin
							mem_ctrl_memorycontroller730 <= verilog_output_f_lhs_array_muxed;
						end
						10'd723: begin
							mem_ctrl_memorycontroller731 <= verilog_output_f_lhs_array_muxed;
						end
						10'd724: begin
							mem_ctrl_memorycontroller732 <= verilog_output_f_lhs_array_muxed;
						end
						10'd725: begin
							mem_ctrl_memorycontroller733 <= verilog_output_f_lhs_array_muxed;
						end
						10'd726: begin
							mem_ctrl_memorycontroller734 <= verilog_output_f_lhs_array_muxed;
						end
						10'd727: begin
							mem_ctrl_memorycontroller735 <= verilog_output_f_lhs_array_muxed;
						end
						10'd728: begin
							mem_ctrl_memorycontroller736 <= verilog_output_f_lhs_array_muxed;
						end
						10'd729: begin
							mem_ctrl_memorycontroller737 <= verilog_output_f_lhs_array_muxed;
						end
						10'd730: begin
							mem_ctrl_memorycontroller738 <= verilog_output_f_lhs_array_muxed;
						end
						10'd731: begin
							mem_ctrl_memorycontroller739 <= verilog_output_f_lhs_array_muxed;
						end
						10'd732: begin
							mem_ctrl_memorycontroller740 <= verilog_output_f_lhs_array_muxed;
						end
						10'd733: begin
							mem_ctrl_memorycontroller741 <= verilog_output_f_lhs_array_muxed;
						end
						10'd734: begin
							mem_ctrl_memorycontroller742 <= verilog_output_f_lhs_array_muxed;
						end
						10'd735: begin
							mem_ctrl_memorycontroller743 <= verilog_output_f_lhs_array_muxed;
						end
						10'd736: begin
							mem_ctrl_memorycontroller744 <= verilog_output_f_lhs_array_muxed;
						end
						10'd737: begin
							mem_ctrl_memorycontroller745 <= verilog_output_f_lhs_array_muxed;
						end
						10'd738: begin
							mem_ctrl_memorycontroller746 <= verilog_output_f_lhs_array_muxed;
						end
						10'd739: begin
							mem_ctrl_memorycontroller747 <= verilog_output_f_lhs_array_muxed;
						end
						10'd740: begin
							mem_ctrl_memorycontroller748 <= verilog_output_f_lhs_array_muxed;
						end
						10'd741: begin
							mem_ctrl_memorycontroller749 <= verilog_output_f_lhs_array_muxed;
						end
						10'd742: begin
							mem_ctrl_memorycontroller750 <= verilog_output_f_lhs_array_muxed;
						end
						10'd743: begin
							mem_ctrl_memorycontroller751 <= verilog_output_f_lhs_array_muxed;
						end
						10'd744: begin
							mem_ctrl_memorycontroller752 <= verilog_output_f_lhs_array_muxed;
						end
						10'd745: begin
							mem_ctrl_memorycontroller753 <= verilog_output_f_lhs_array_muxed;
						end
						10'd746: begin
							mem_ctrl_memorycontroller754 <= verilog_output_f_lhs_array_muxed;
						end
						10'd747: begin
							mem_ctrl_memorycontroller755 <= verilog_output_f_lhs_array_muxed;
						end
						10'd748: begin
							mem_ctrl_memorycontroller756 <= verilog_output_f_lhs_array_muxed;
						end
						10'd749: begin
							mem_ctrl_memorycontroller757 <= verilog_output_f_lhs_array_muxed;
						end
						10'd750: begin
							mem_ctrl_memorycontroller758 <= verilog_output_f_lhs_array_muxed;
						end
						10'd751: begin
							mem_ctrl_memorycontroller759 <= verilog_output_f_lhs_array_muxed;
						end
						10'd752: begin
							mem_ctrl_memorycontroller760 <= verilog_output_f_lhs_array_muxed;
						end
						10'd753: begin
							mem_ctrl_memorycontroller761 <= verilog_output_f_lhs_array_muxed;
						end
						10'd754: begin
							mem_ctrl_memorycontroller762 <= verilog_output_f_lhs_array_muxed;
						end
						10'd755: begin
							mem_ctrl_memorycontroller763 <= verilog_output_f_lhs_array_muxed;
						end
						10'd756: begin
							mem_ctrl_memorycontroller764 <= verilog_output_f_lhs_array_muxed;
						end
						10'd757: begin
							mem_ctrl_memorycontroller765 <= verilog_output_f_lhs_array_muxed;
						end
						10'd758: begin
							mem_ctrl_memorycontroller766 <= verilog_output_f_lhs_array_muxed;
						end
						10'd759: begin
							mem_ctrl_memorycontroller767 <= verilog_output_f_lhs_array_muxed;
						end
						10'd760: begin
							mem_ctrl_memorycontroller768 <= verilog_output_f_lhs_array_muxed;
						end
						10'd761: begin
							mem_ctrl_memorycontroller769 <= verilog_output_f_lhs_array_muxed;
						end
						10'd762: begin
							mem_ctrl_memorycontroller770 <= verilog_output_f_lhs_array_muxed;
						end
						10'd763: begin
							mem_ctrl_memorycontroller771 <= verilog_output_f_lhs_array_muxed;
						end
						10'd764: begin
							mem_ctrl_memorycontroller772 <= verilog_output_f_lhs_array_muxed;
						end
						10'd765: begin
							mem_ctrl_memorycontroller773 <= verilog_output_f_lhs_array_muxed;
						end
						10'd766: begin
							mem_ctrl_memorycontroller774 <= verilog_output_f_lhs_array_muxed;
						end
						10'd767: begin
							mem_ctrl_memorycontroller775 <= verilog_output_f_lhs_array_muxed;
						end
						10'd768: begin
							mem_ctrl_memorycontroller776 <= verilog_output_f_lhs_array_muxed;
						end
						10'd769: begin
							mem_ctrl_memorycontroller777 <= verilog_output_f_lhs_array_muxed;
						end
						10'd770: begin
							mem_ctrl_memorycontroller778 <= verilog_output_f_lhs_array_muxed;
						end
						10'd771: begin
							mem_ctrl_memorycontroller779 <= verilog_output_f_lhs_array_muxed;
						end
						10'd772: begin
							mem_ctrl_memorycontroller780 <= verilog_output_f_lhs_array_muxed;
						end
						10'd773: begin
							mem_ctrl_memorycontroller781 <= verilog_output_f_lhs_array_muxed;
						end
						10'd774: begin
							mem_ctrl_memorycontroller782 <= verilog_output_f_lhs_array_muxed;
						end
						10'd775: begin
							mem_ctrl_memorycontroller783 <= verilog_output_f_lhs_array_muxed;
						end
						10'd776: begin
							mem_ctrl_memorycontroller784 <= verilog_output_f_lhs_array_muxed;
						end
						10'd777: begin
							mem_ctrl_memorycontroller785 <= verilog_output_f_lhs_array_muxed;
						end
						10'd778: begin
							mem_ctrl_memorycontroller786 <= verilog_output_f_lhs_array_muxed;
						end
						10'd779: begin
							mem_ctrl_memorycontroller787 <= verilog_output_f_lhs_array_muxed;
						end
						10'd780: begin
							mem_ctrl_memorycontroller788 <= verilog_output_f_lhs_array_muxed;
						end
						10'd781: begin
							mem_ctrl_memorycontroller789 <= verilog_output_f_lhs_array_muxed;
						end
						10'd782: begin
							mem_ctrl_memorycontroller790 <= verilog_output_f_lhs_array_muxed;
						end
						10'd783: begin
							mem_ctrl_memorycontroller791 <= verilog_output_f_lhs_array_muxed;
						end
						10'd784: begin
							mem_ctrl_memorycontroller792 <= verilog_output_f_lhs_array_muxed;
						end
						10'd785: begin
							mem_ctrl_memorycontroller793 <= verilog_output_f_lhs_array_muxed;
						end
						10'd786: begin
							mem_ctrl_memorycontroller794 <= verilog_output_f_lhs_array_muxed;
						end
						10'd787: begin
							mem_ctrl_memorycontroller795 <= verilog_output_f_lhs_array_muxed;
						end
						10'd788: begin
							mem_ctrl_memorycontroller796 <= verilog_output_f_lhs_array_muxed;
						end
						10'd789: begin
							mem_ctrl_memorycontroller797 <= verilog_output_f_lhs_array_muxed;
						end
						10'd790: begin
							mem_ctrl_memorycontroller798 <= verilog_output_f_lhs_array_muxed;
						end
						10'd791: begin
							mem_ctrl_memorycontroller799 <= verilog_output_f_lhs_array_muxed;
						end
						10'd792: begin
							mem_ctrl_memorycontroller800 <= verilog_output_f_lhs_array_muxed;
						end
						10'd793: begin
							mem_ctrl_memorycontroller801 <= verilog_output_f_lhs_array_muxed;
						end
						10'd794: begin
							mem_ctrl_memorycontroller802 <= verilog_output_f_lhs_array_muxed;
						end
						10'd795: begin
							mem_ctrl_memorycontroller803 <= verilog_output_f_lhs_array_muxed;
						end
						10'd796: begin
							mem_ctrl_memorycontroller804 <= verilog_output_f_lhs_array_muxed;
						end
						10'd797: begin
							mem_ctrl_memorycontroller805 <= verilog_output_f_lhs_array_muxed;
						end
						10'd798: begin
							mem_ctrl_memorycontroller806 <= verilog_output_f_lhs_array_muxed;
						end
						10'd799: begin
							mem_ctrl_memorycontroller807 <= verilog_output_f_lhs_array_muxed;
						end
						10'd800: begin
							mem_ctrl_memorycontroller808 <= verilog_output_f_lhs_array_muxed;
						end
						10'd801: begin
							mem_ctrl_memorycontroller809 <= verilog_output_f_lhs_array_muxed;
						end
						10'd802: begin
							mem_ctrl_memorycontroller810 <= verilog_output_f_lhs_array_muxed;
						end
						10'd803: begin
							mem_ctrl_memorycontroller811 <= verilog_output_f_lhs_array_muxed;
						end
						10'd804: begin
							mem_ctrl_memorycontroller812 <= verilog_output_f_lhs_array_muxed;
						end
						10'd805: begin
							mem_ctrl_memorycontroller813 <= verilog_output_f_lhs_array_muxed;
						end
						10'd806: begin
							mem_ctrl_memorycontroller814 <= verilog_output_f_lhs_array_muxed;
						end
						10'd807: begin
							mem_ctrl_memorycontroller815 <= verilog_output_f_lhs_array_muxed;
						end
						10'd808: begin
							mem_ctrl_memorycontroller816 <= verilog_output_f_lhs_array_muxed;
						end
						10'd809: begin
							mem_ctrl_memorycontroller817 <= verilog_output_f_lhs_array_muxed;
						end
						10'd810: begin
							mem_ctrl_memorycontroller818 <= verilog_output_f_lhs_array_muxed;
						end
						10'd811: begin
							mem_ctrl_memorycontroller819 <= verilog_output_f_lhs_array_muxed;
						end
						10'd812: begin
							mem_ctrl_memorycontroller820 <= verilog_output_f_lhs_array_muxed;
						end
						10'd813: begin
							mem_ctrl_memorycontroller821 <= verilog_output_f_lhs_array_muxed;
						end
						10'd814: begin
							mem_ctrl_memorycontroller822 <= verilog_output_f_lhs_array_muxed;
						end
						10'd815: begin
							mem_ctrl_memorycontroller823 <= verilog_output_f_lhs_array_muxed;
						end
						10'd816: begin
							mem_ctrl_memorycontroller824 <= verilog_output_f_lhs_array_muxed;
						end
						10'd817: begin
							mem_ctrl_memorycontroller825 <= verilog_output_f_lhs_array_muxed;
						end
						10'd818: begin
							mem_ctrl_memorycontroller826 <= verilog_output_f_lhs_array_muxed;
						end
						10'd819: begin
							mem_ctrl_memorycontroller827 <= verilog_output_f_lhs_array_muxed;
						end
						10'd820: begin
							mem_ctrl_memorycontroller828 <= verilog_output_f_lhs_array_muxed;
						end
						10'd821: begin
							mem_ctrl_memorycontroller829 <= verilog_output_f_lhs_array_muxed;
						end
						10'd822: begin
							mem_ctrl_memorycontroller830 <= verilog_output_f_lhs_array_muxed;
						end
						10'd823: begin
							mem_ctrl_memorycontroller831 <= verilog_output_f_lhs_array_muxed;
						end
						10'd824: begin
							mem_ctrl_memorycontroller832 <= verilog_output_f_lhs_array_muxed;
						end
						10'd825: begin
							mem_ctrl_memorycontroller833 <= verilog_output_f_lhs_array_muxed;
						end
						10'd826: begin
							mem_ctrl_memorycontroller834 <= verilog_output_f_lhs_array_muxed;
						end
						10'd827: begin
							mem_ctrl_memorycontroller835 <= verilog_output_f_lhs_array_muxed;
						end
						10'd828: begin
							mem_ctrl_memorycontroller836 <= verilog_output_f_lhs_array_muxed;
						end
						10'd829: begin
							mem_ctrl_memorycontroller837 <= verilog_output_f_lhs_array_muxed;
						end
						10'd830: begin
							mem_ctrl_memorycontroller838 <= verilog_output_f_lhs_array_muxed;
						end
						10'd831: begin
							mem_ctrl_memorycontroller839 <= verilog_output_f_lhs_array_muxed;
						end
						10'd832: begin
							mem_ctrl_memorycontroller840 <= verilog_output_f_lhs_array_muxed;
						end
						10'd833: begin
							mem_ctrl_memorycontroller841 <= verilog_output_f_lhs_array_muxed;
						end
						10'd834: begin
							mem_ctrl_memorycontroller842 <= verilog_output_f_lhs_array_muxed;
						end
						10'd835: begin
							mem_ctrl_memorycontroller843 <= verilog_output_f_lhs_array_muxed;
						end
						10'd836: begin
							mem_ctrl_memorycontroller844 <= verilog_output_f_lhs_array_muxed;
						end
						10'd837: begin
							mem_ctrl_memorycontroller845 <= verilog_output_f_lhs_array_muxed;
						end
						10'd838: begin
							mem_ctrl_memorycontroller846 <= verilog_output_f_lhs_array_muxed;
						end
						10'd839: begin
							mem_ctrl_memorycontroller847 <= verilog_output_f_lhs_array_muxed;
						end
						10'd840: begin
							mem_ctrl_memorycontroller848 <= verilog_output_f_lhs_array_muxed;
						end
						10'd841: begin
							mem_ctrl_memorycontroller849 <= verilog_output_f_lhs_array_muxed;
						end
						10'd842: begin
							mem_ctrl_memorycontroller850 <= verilog_output_f_lhs_array_muxed;
						end
						10'd843: begin
							mem_ctrl_memorycontroller851 <= verilog_output_f_lhs_array_muxed;
						end
						10'd844: begin
							mem_ctrl_memorycontroller852 <= verilog_output_f_lhs_array_muxed;
						end
						10'd845: begin
							mem_ctrl_memorycontroller853 <= verilog_output_f_lhs_array_muxed;
						end
						10'd846: begin
							mem_ctrl_memorycontroller854 <= verilog_output_f_lhs_array_muxed;
						end
						10'd847: begin
							mem_ctrl_memorycontroller855 <= verilog_output_f_lhs_array_muxed;
						end
						10'd848: begin
							mem_ctrl_memorycontroller856 <= verilog_output_f_lhs_array_muxed;
						end
						10'd849: begin
							mem_ctrl_memorycontroller857 <= verilog_output_f_lhs_array_muxed;
						end
						10'd850: begin
							mem_ctrl_memorycontroller858 <= verilog_output_f_lhs_array_muxed;
						end
						10'd851: begin
							mem_ctrl_memorycontroller859 <= verilog_output_f_lhs_array_muxed;
						end
						10'd852: begin
							mem_ctrl_memorycontroller860 <= verilog_output_f_lhs_array_muxed;
						end
						10'd853: begin
							mem_ctrl_memorycontroller861 <= verilog_output_f_lhs_array_muxed;
						end
						10'd854: begin
							mem_ctrl_memorycontroller862 <= verilog_output_f_lhs_array_muxed;
						end
						10'd855: begin
							mem_ctrl_memorycontroller863 <= verilog_output_f_lhs_array_muxed;
						end
						10'd856: begin
							mem_ctrl_memorycontroller864 <= verilog_output_f_lhs_array_muxed;
						end
						10'd857: begin
							mem_ctrl_memorycontroller865 <= verilog_output_f_lhs_array_muxed;
						end
						10'd858: begin
							mem_ctrl_memorycontroller866 <= verilog_output_f_lhs_array_muxed;
						end
						10'd859: begin
							mem_ctrl_memorycontroller867 <= verilog_output_f_lhs_array_muxed;
						end
						10'd860: begin
							mem_ctrl_memorycontroller868 <= verilog_output_f_lhs_array_muxed;
						end
						10'd861: begin
							mem_ctrl_memorycontroller869 <= verilog_output_f_lhs_array_muxed;
						end
						10'd862: begin
							mem_ctrl_memorycontroller870 <= verilog_output_f_lhs_array_muxed;
						end
						10'd863: begin
							mem_ctrl_memorycontroller871 <= verilog_output_f_lhs_array_muxed;
						end
						10'd864: begin
							mem_ctrl_memorycontroller872 <= verilog_output_f_lhs_array_muxed;
						end
						10'd865: begin
							mem_ctrl_memorycontroller873 <= verilog_output_f_lhs_array_muxed;
						end
						10'd866: begin
							mem_ctrl_memorycontroller874 <= verilog_output_f_lhs_array_muxed;
						end
						10'd867: begin
							mem_ctrl_memorycontroller875 <= verilog_output_f_lhs_array_muxed;
						end
						10'd868: begin
							mem_ctrl_memorycontroller876 <= verilog_output_f_lhs_array_muxed;
						end
						10'd869: begin
							mem_ctrl_memorycontroller877 <= verilog_output_f_lhs_array_muxed;
						end
						10'd870: begin
							mem_ctrl_memorycontroller878 <= verilog_output_f_lhs_array_muxed;
						end
						10'd871: begin
							mem_ctrl_memorycontroller879 <= verilog_output_f_lhs_array_muxed;
						end
						10'd872: begin
							mem_ctrl_memorycontroller880 <= verilog_output_f_lhs_array_muxed;
						end
						10'd873: begin
							mem_ctrl_memorycontroller881 <= verilog_output_f_lhs_array_muxed;
						end
						10'd874: begin
							mem_ctrl_memorycontroller882 <= verilog_output_f_lhs_array_muxed;
						end
						10'd875: begin
							mem_ctrl_memorycontroller883 <= verilog_output_f_lhs_array_muxed;
						end
						10'd876: begin
							mem_ctrl_memorycontroller884 <= verilog_output_f_lhs_array_muxed;
						end
						10'd877: begin
							mem_ctrl_memorycontroller885 <= verilog_output_f_lhs_array_muxed;
						end
						10'd878: begin
							mem_ctrl_memorycontroller886 <= verilog_output_f_lhs_array_muxed;
						end
						10'd879: begin
							mem_ctrl_memorycontroller887 <= verilog_output_f_lhs_array_muxed;
						end
						10'd880: begin
							mem_ctrl_memorycontroller888 <= verilog_output_f_lhs_array_muxed;
						end
						10'd881: begin
							mem_ctrl_memorycontroller889 <= verilog_output_f_lhs_array_muxed;
						end
						10'd882: begin
							mem_ctrl_memorycontroller890 <= verilog_output_f_lhs_array_muxed;
						end
						10'd883: begin
							mem_ctrl_memorycontroller891 <= verilog_output_f_lhs_array_muxed;
						end
						10'd884: begin
							mem_ctrl_memorycontroller892 <= verilog_output_f_lhs_array_muxed;
						end
						10'd885: begin
							mem_ctrl_memorycontroller893 <= verilog_output_f_lhs_array_muxed;
						end
						10'd886: begin
							mem_ctrl_memorycontroller894 <= verilog_output_f_lhs_array_muxed;
						end
						10'd887: begin
							mem_ctrl_memorycontroller895 <= verilog_output_f_lhs_array_muxed;
						end
						10'd888: begin
							mem_ctrl_memorycontroller896 <= verilog_output_f_lhs_array_muxed;
						end
						10'd889: begin
							mem_ctrl_memorycontroller897 <= verilog_output_f_lhs_array_muxed;
						end
						10'd890: begin
							mem_ctrl_memorycontroller898 <= verilog_output_f_lhs_array_muxed;
						end
						10'd891: begin
							mem_ctrl_memorycontroller899 <= verilog_output_f_lhs_array_muxed;
						end
						10'd892: begin
							mem_ctrl_memorycontroller900 <= verilog_output_f_lhs_array_muxed;
						end
						10'd893: begin
							mem_ctrl_memorycontroller901 <= verilog_output_f_lhs_array_muxed;
						end
						10'd894: begin
							mem_ctrl_memorycontroller902 <= verilog_output_f_lhs_array_muxed;
						end
						10'd895: begin
							mem_ctrl_memorycontroller903 <= verilog_output_f_lhs_array_muxed;
						end
						10'd896: begin
							mem_ctrl_memorycontroller904 <= verilog_output_f_lhs_array_muxed;
						end
						10'd897: begin
							mem_ctrl_memorycontroller905 <= verilog_output_f_lhs_array_muxed;
						end
						10'd898: begin
							mem_ctrl_memorycontroller906 <= verilog_output_f_lhs_array_muxed;
						end
						10'd899: begin
							mem_ctrl_memorycontroller907 <= verilog_output_f_lhs_array_muxed;
						end
						10'd900: begin
							mem_ctrl_memorycontroller908 <= verilog_output_f_lhs_array_muxed;
						end
						10'd901: begin
							mem_ctrl_memorycontroller909 <= verilog_output_f_lhs_array_muxed;
						end
						10'd902: begin
							mem_ctrl_memorycontroller910 <= verilog_output_f_lhs_array_muxed;
						end
						10'd903: begin
							mem_ctrl_memorycontroller911 <= verilog_output_f_lhs_array_muxed;
						end
						10'd904: begin
							mem_ctrl_memorycontroller912 <= verilog_output_f_lhs_array_muxed;
						end
						10'd905: begin
							mem_ctrl_memorycontroller913 <= verilog_output_f_lhs_array_muxed;
						end
						10'd906: begin
							mem_ctrl_memorycontroller914 <= verilog_output_f_lhs_array_muxed;
						end
						10'd907: begin
							mem_ctrl_memorycontroller915 <= verilog_output_f_lhs_array_muxed;
						end
						10'd908: begin
							mem_ctrl_memorycontroller916 <= verilog_output_f_lhs_array_muxed;
						end
						10'd909: begin
							mem_ctrl_memorycontroller917 <= verilog_output_f_lhs_array_muxed;
						end
						10'd910: begin
							mem_ctrl_memorycontroller918 <= verilog_output_f_lhs_array_muxed;
						end
						10'd911: begin
							mem_ctrl_memorycontroller919 <= verilog_output_f_lhs_array_muxed;
						end
						10'd912: begin
							mem_ctrl_memorycontroller920 <= verilog_output_f_lhs_array_muxed;
						end
						10'd913: begin
							mem_ctrl_memorycontroller921 <= verilog_output_f_lhs_array_muxed;
						end
						10'd914: begin
							mem_ctrl_memorycontroller922 <= verilog_output_f_lhs_array_muxed;
						end
						10'd915: begin
							mem_ctrl_memorycontroller923 <= verilog_output_f_lhs_array_muxed;
						end
						10'd916: begin
							mem_ctrl_memorycontroller924 <= verilog_output_f_lhs_array_muxed;
						end
						10'd917: begin
							mem_ctrl_memorycontroller925 <= verilog_output_f_lhs_array_muxed;
						end
						10'd918: begin
							mem_ctrl_memorycontroller926 <= verilog_output_f_lhs_array_muxed;
						end
						10'd919: begin
							mem_ctrl_memorycontroller927 <= verilog_output_f_lhs_array_muxed;
						end
						10'd920: begin
							mem_ctrl_memorycontroller928 <= verilog_output_f_lhs_array_muxed;
						end
						10'd921: begin
							mem_ctrl_memorycontroller929 <= verilog_output_f_lhs_array_muxed;
						end
						10'd922: begin
							mem_ctrl_memorycontroller930 <= verilog_output_f_lhs_array_muxed;
						end
						10'd923: begin
							mem_ctrl_memorycontroller931 <= verilog_output_f_lhs_array_muxed;
						end
						10'd924: begin
							mem_ctrl_memorycontroller932 <= verilog_output_f_lhs_array_muxed;
						end
						10'd925: begin
							mem_ctrl_memorycontroller933 <= verilog_output_f_lhs_array_muxed;
						end
						10'd926: begin
							mem_ctrl_memorycontroller934 <= verilog_output_f_lhs_array_muxed;
						end
						10'd927: begin
							mem_ctrl_memorycontroller935 <= verilog_output_f_lhs_array_muxed;
						end
						10'd928: begin
							mem_ctrl_memorycontroller936 <= verilog_output_f_lhs_array_muxed;
						end
						10'd929: begin
							mem_ctrl_memorycontroller937 <= verilog_output_f_lhs_array_muxed;
						end
						10'd930: begin
							mem_ctrl_memorycontroller938 <= verilog_output_f_lhs_array_muxed;
						end
						10'd931: begin
							mem_ctrl_memorycontroller939 <= verilog_output_f_lhs_array_muxed;
						end
						10'd932: begin
							mem_ctrl_memorycontroller940 <= verilog_output_f_lhs_array_muxed;
						end
						10'd933: begin
							mem_ctrl_memorycontroller941 <= verilog_output_f_lhs_array_muxed;
						end
						10'd934: begin
							mem_ctrl_memorycontroller942 <= verilog_output_f_lhs_array_muxed;
						end
						10'd935: begin
							mem_ctrl_memorycontroller943 <= verilog_output_f_lhs_array_muxed;
						end
						10'd936: begin
							mem_ctrl_memorycontroller944 <= verilog_output_f_lhs_array_muxed;
						end
						10'd937: begin
							mem_ctrl_memorycontroller945 <= verilog_output_f_lhs_array_muxed;
						end
						10'd938: begin
							mem_ctrl_memorycontroller946 <= verilog_output_f_lhs_array_muxed;
						end
						10'd939: begin
							mem_ctrl_memorycontroller947 <= verilog_output_f_lhs_array_muxed;
						end
						10'd940: begin
							mem_ctrl_memorycontroller948 <= verilog_output_f_lhs_array_muxed;
						end
						10'd941: begin
							mem_ctrl_memorycontroller949 <= verilog_output_f_lhs_array_muxed;
						end
						10'd942: begin
							mem_ctrl_memorycontroller950 <= verilog_output_f_lhs_array_muxed;
						end
						10'd943: begin
							mem_ctrl_memorycontroller951 <= verilog_output_f_lhs_array_muxed;
						end
						10'd944: begin
							mem_ctrl_memorycontroller952 <= verilog_output_f_lhs_array_muxed;
						end
						10'd945: begin
							mem_ctrl_memorycontroller953 <= verilog_output_f_lhs_array_muxed;
						end
						10'd946: begin
							mem_ctrl_memorycontroller954 <= verilog_output_f_lhs_array_muxed;
						end
						10'd947: begin
							mem_ctrl_memorycontroller955 <= verilog_output_f_lhs_array_muxed;
						end
						10'd948: begin
							mem_ctrl_memorycontroller956 <= verilog_output_f_lhs_array_muxed;
						end
						10'd949: begin
							mem_ctrl_memorycontroller957 <= verilog_output_f_lhs_array_muxed;
						end
						10'd950: begin
							mem_ctrl_memorycontroller958 <= verilog_output_f_lhs_array_muxed;
						end
						10'd951: begin
							mem_ctrl_memorycontroller959 <= verilog_output_f_lhs_array_muxed;
						end
						10'd952: begin
							mem_ctrl_memorycontroller960 <= verilog_output_f_lhs_array_muxed;
						end
						10'd953: begin
							mem_ctrl_memorycontroller961 <= verilog_output_f_lhs_array_muxed;
						end
						10'd954: begin
							mem_ctrl_memorycontroller962 <= verilog_output_f_lhs_array_muxed;
						end
						10'd955: begin
							mem_ctrl_memorycontroller963 <= verilog_output_f_lhs_array_muxed;
						end
						10'd956: begin
							mem_ctrl_memorycontroller964 <= verilog_output_f_lhs_array_muxed;
						end
						10'd957: begin
							mem_ctrl_memorycontroller965 <= verilog_output_f_lhs_array_muxed;
						end
						10'd958: begin
							mem_ctrl_memorycontroller966 <= verilog_output_f_lhs_array_muxed;
						end
						10'd959: begin
							mem_ctrl_memorycontroller967 <= verilog_output_f_lhs_array_muxed;
						end
						10'd960: begin
							mem_ctrl_memorycontroller968 <= verilog_output_f_lhs_array_muxed;
						end
						10'd961: begin
							mem_ctrl_memorycontroller969 <= verilog_output_f_lhs_array_muxed;
						end
						10'd962: begin
							mem_ctrl_memorycontroller970 <= verilog_output_f_lhs_array_muxed;
						end
						10'd963: begin
							mem_ctrl_memorycontroller971 <= verilog_output_f_lhs_array_muxed;
						end
						10'd964: begin
							mem_ctrl_memorycontroller972 <= verilog_output_f_lhs_array_muxed;
						end
						10'd965: begin
							mem_ctrl_memorycontroller973 <= verilog_output_f_lhs_array_muxed;
						end
						10'd966: begin
							mem_ctrl_memorycontroller974 <= verilog_output_f_lhs_array_muxed;
						end
						10'd967: begin
							mem_ctrl_memorycontroller975 <= verilog_output_f_lhs_array_muxed;
						end
						10'd968: begin
							mem_ctrl_memorycontroller976 <= verilog_output_f_lhs_array_muxed;
						end
						10'd969: begin
							mem_ctrl_memorycontroller977 <= verilog_output_f_lhs_array_muxed;
						end
						10'd970: begin
							mem_ctrl_memorycontroller978 <= verilog_output_f_lhs_array_muxed;
						end
						10'd971: begin
							mem_ctrl_memorycontroller979 <= verilog_output_f_lhs_array_muxed;
						end
						10'd972: begin
							mem_ctrl_memorycontroller980 <= verilog_output_f_lhs_array_muxed;
						end
						10'd973: begin
							mem_ctrl_memorycontroller981 <= verilog_output_f_lhs_array_muxed;
						end
						10'd974: begin
							mem_ctrl_memorycontroller982 <= verilog_output_f_lhs_array_muxed;
						end
						10'd975: begin
							mem_ctrl_memorycontroller983 <= verilog_output_f_lhs_array_muxed;
						end
						10'd976: begin
							mem_ctrl_memorycontroller984 <= verilog_output_f_lhs_array_muxed;
						end
						10'd977: begin
							mem_ctrl_memorycontroller985 <= verilog_output_f_lhs_array_muxed;
						end
						10'd978: begin
							mem_ctrl_memorycontroller986 <= verilog_output_f_lhs_array_muxed;
						end
						10'd979: begin
							mem_ctrl_memorycontroller987 <= verilog_output_f_lhs_array_muxed;
						end
						10'd980: begin
							mem_ctrl_memorycontroller988 <= verilog_output_f_lhs_array_muxed;
						end
						10'd981: begin
							mem_ctrl_memorycontroller989 <= verilog_output_f_lhs_array_muxed;
						end
						10'd982: begin
							mem_ctrl_memorycontroller990 <= verilog_output_f_lhs_array_muxed;
						end
						10'd983: begin
							mem_ctrl_memorycontroller991 <= verilog_output_f_lhs_array_muxed;
						end
						10'd984: begin
							mem_ctrl_memorycontroller992 <= verilog_output_f_lhs_array_muxed;
						end
						10'd985: begin
							mem_ctrl_memorycontroller993 <= verilog_output_f_lhs_array_muxed;
						end
						10'd986: begin
							mem_ctrl_memorycontroller994 <= verilog_output_f_lhs_array_muxed;
						end
						10'd987: begin
							mem_ctrl_memorycontroller995 <= verilog_output_f_lhs_array_muxed;
						end
						10'd988: begin
							mem_ctrl_memorycontroller996 <= verilog_output_f_lhs_array_muxed;
						end
						10'd989: begin
							mem_ctrl_memorycontroller997 <= verilog_output_f_lhs_array_muxed;
						end
						10'd990: begin
							mem_ctrl_memorycontroller998 <= verilog_output_f_lhs_array_muxed;
						end
						10'd991: begin
							mem_ctrl_memorycontroller999 <= verilog_output_f_lhs_array_muxed;
						end
						10'd992: begin
							mem_ctrl_memorycontroller1000 <= verilog_output_f_lhs_array_muxed;
						end
						10'd993: begin
							mem_ctrl_memorycontroller1001 <= verilog_output_f_lhs_array_muxed;
						end
						10'd994: begin
							mem_ctrl_memorycontroller1002 <= verilog_output_f_lhs_array_muxed;
						end
						10'd995: begin
							mem_ctrl_memorycontroller1003 <= verilog_output_f_lhs_array_muxed;
						end
						10'd996: begin
							mem_ctrl_memorycontroller1004 <= verilog_output_f_lhs_array_muxed;
						end
						10'd997: begin
							mem_ctrl_memorycontroller1005 <= verilog_output_f_lhs_array_muxed;
						end
						10'd998: begin
							mem_ctrl_memorycontroller1006 <= verilog_output_f_lhs_array_muxed;
						end
						10'd999: begin
							mem_ctrl_memorycontroller1007 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1000: begin
							mem_ctrl_memorycontroller1008 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1001: begin
							mem_ctrl_memorycontroller1009 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1002: begin
							mem_ctrl_memorycontroller1010 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1003: begin
							mem_ctrl_memorycontroller1011 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1004: begin
							mem_ctrl_memorycontroller1012 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1005: begin
							mem_ctrl_memorycontroller1013 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1006: begin
							mem_ctrl_memorycontroller1014 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1007: begin
							mem_ctrl_memorycontroller1015 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1008: begin
							mem_ctrl_memorycontroller1016 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1009: begin
							mem_ctrl_memorycontroller1017 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1010: begin
							mem_ctrl_memorycontroller1018 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1011: begin
							mem_ctrl_memorycontroller1019 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1012: begin
							mem_ctrl_memorycontroller1020 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1013: begin
							mem_ctrl_memorycontroller1021 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1014: begin
							mem_ctrl_memorycontroller1022 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1015: begin
							mem_ctrl_memorycontroller1023 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1016: begin
							mem_ctrl_memorycontroller1024 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1017: begin
							mem_ctrl_memorycontroller1025 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1018: begin
							mem_ctrl_memorycontroller1026 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1019: begin
							mem_ctrl_memorycontroller1027 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1020: begin
							mem_ctrl_memorycontroller1028 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1021: begin
							mem_ctrl_memorycontroller1029 <= verilog_output_f_lhs_array_muxed;
						end
						10'd1022: begin
							mem_ctrl_memorycontroller1030 <= verilog_output_f_lhs_array_muxed;
						end
						default: begin
							mem_ctrl_memorycontroller1031 <= verilog_output_f_lhs_array_muxed;
						end
					endcase
				end
			end
		end
	end
	if (sys_rst) begin
		data_out <= 64'd0;
		ready <= 1'd0;
		mem_ctrl_cmd_decoded <= 4'd0;
		mem_ctrl_address <= 32'd0;
		mem_ctrl_timer <= 32'd0;
		mem_ctrl_state <= 2'd0;
		mem_ctrl_memorycontroller0 <= 64'd0;
		mem_ctrl_memorycontroller1 <= 64'd0;
		mem_ctrl_memorycontroller2 <= 64'd0;
		mem_ctrl_memorycontroller3 <= 64'd0;
		mem_ctrl_memorycontroller4 <= 64'd0;
		mem_ctrl_memorycontroller5 <= 64'd0;
		mem_ctrl_memorycontroller6 <= 64'd0;
		mem_ctrl_memorycontroller7 <= 64'd0;
		mem_ctrl_buffer_index <= 3'd0;
		mem_ctrl_power_state <= 2'd0;
		mem_ctrl_memorycontroller8 <= 64'd0;
		mem_ctrl_memorycontroller9 <= 64'd0;
		mem_ctrl_memorycontroller10 <= 64'd0;
		mem_ctrl_memorycontroller11 <= 64'd0;
		mem_ctrl_memorycontroller12 <= 64'd0;
		mem_ctrl_memorycontroller13 <= 64'd0;
		mem_ctrl_memorycontroller14 <= 64'd0;
		mem_ctrl_memorycontroller15 <= 64'd0;
		mem_ctrl_memorycontroller16 <= 64'd0;
		mem_ctrl_memorycontroller17 <= 64'd0;
		mem_ctrl_memorycontroller18 <= 64'd0;
		mem_ctrl_memorycontroller19 <= 64'd0;
		mem_ctrl_memorycontroller20 <= 64'd0;
		mem_ctrl_memorycontroller21 <= 64'd0;
		mem_ctrl_memorycontroller22 <= 64'd0;
		mem_ctrl_memorycontroller23 <= 64'd0;
		mem_ctrl_memorycontroller24 <= 64'd0;
		mem_ctrl_memorycontroller25 <= 64'd0;
		mem_ctrl_memorycontroller26 <= 64'd0;
		mem_ctrl_memorycontroller27 <= 64'd0;
		mem_ctrl_memorycontroller28 <= 64'd0;
		mem_ctrl_memorycontroller29 <= 64'd0;
		mem_ctrl_memorycontroller30 <= 64'd0;
		mem_ctrl_memorycontroller31 <= 64'd0;
		mem_ctrl_memorycontroller32 <= 64'd0;
		mem_ctrl_memorycontroller33 <= 64'd0;
		mem_ctrl_memorycontroller34 <= 64'd0;
		mem_ctrl_memorycontroller35 <= 64'd0;
		mem_ctrl_memorycontroller36 <= 64'd0;
		mem_ctrl_memorycontroller37 <= 64'd0;
		mem_ctrl_memorycontroller38 <= 64'd0;
		mem_ctrl_memorycontroller39 <= 64'd0;
		mem_ctrl_memorycontroller40 <= 64'd0;
		mem_ctrl_memorycontroller41 <= 64'd0;
		mem_ctrl_memorycontroller42 <= 64'd0;
		mem_ctrl_memorycontroller43 <= 64'd0;
		mem_ctrl_memorycontroller44 <= 64'd0;
		mem_ctrl_memorycontroller45 <= 64'd0;
		mem_ctrl_memorycontroller46 <= 64'd0;
		mem_ctrl_memorycontroller47 <= 64'd0;
		mem_ctrl_memorycontroller48 <= 64'd0;
		mem_ctrl_memorycontroller49 <= 64'd0;
		mem_ctrl_memorycontroller50 <= 64'd0;
		mem_ctrl_memorycontroller51 <= 64'd0;
		mem_ctrl_memorycontroller52 <= 64'd0;
		mem_ctrl_memorycontroller53 <= 64'd0;
		mem_ctrl_memorycontroller54 <= 64'd0;
		mem_ctrl_memorycontroller55 <= 64'd0;
		mem_ctrl_memorycontroller56 <= 64'd0;
		mem_ctrl_memorycontroller57 <= 64'd0;
		mem_ctrl_memorycontroller58 <= 64'd0;
		mem_ctrl_memorycontroller59 <= 64'd0;
		mem_ctrl_memorycontroller60 <= 64'd0;
		mem_ctrl_memorycontroller61 <= 64'd0;
		mem_ctrl_memorycontroller62 <= 64'd0;
		mem_ctrl_memorycontroller63 <= 64'd0;
		mem_ctrl_memorycontroller64 <= 64'd0;
		mem_ctrl_memorycontroller65 <= 64'd0;
		mem_ctrl_memorycontroller66 <= 64'd0;
		mem_ctrl_memorycontroller67 <= 64'd0;
		mem_ctrl_memorycontroller68 <= 64'd0;
		mem_ctrl_memorycontroller69 <= 64'd0;
		mem_ctrl_memorycontroller70 <= 64'd0;
		mem_ctrl_memorycontroller71 <= 64'd0;
		mem_ctrl_memorycontroller72 <= 64'd0;
		mem_ctrl_memorycontroller73 <= 64'd0;
		mem_ctrl_memorycontroller74 <= 64'd0;
		mem_ctrl_memorycontroller75 <= 64'd0;
		mem_ctrl_memorycontroller76 <= 64'd0;
		mem_ctrl_memorycontroller77 <= 64'd0;
		mem_ctrl_memorycontroller78 <= 64'd0;
		mem_ctrl_memorycontroller79 <= 64'd0;
		mem_ctrl_memorycontroller80 <= 64'd0;
		mem_ctrl_memorycontroller81 <= 64'd0;
		mem_ctrl_memorycontroller82 <= 64'd0;
		mem_ctrl_memorycontroller83 <= 64'd0;
		mem_ctrl_memorycontroller84 <= 64'd0;
		mem_ctrl_memorycontroller85 <= 64'd0;
		mem_ctrl_memorycontroller86 <= 64'd0;
		mem_ctrl_memorycontroller87 <= 64'd0;
		mem_ctrl_memorycontroller88 <= 64'd0;
		mem_ctrl_memorycontroller89 <= 64'd0;
		mem_ctrl_memorycontroller90 <= 64'd0;
		mem_ctrl_memorycontroller91 <= 64'd0;
		mem_ctrl_memorycontroller92 <= 64'd0;
		mem_ctrl_memorycontroller93 <= 64'd0;
		mem_ctrl_memorycontroller94 <= 64'd0;
		mem_ctrl_memorycontroller95 <= 64'd0;
		mem_ctrl_memorycontroller96 <= 64'd0;
		mem_ctrl_memorycontroller97 <= 64'd0;
		mem_ctrl_memorycontroller98 <= 64'd0;
		mem_ctrl_memorycontroller99 <= 64'd0;
		mem_ctrl_memorycontroller100 <= 64'd0;
		mem_ctrl_memorycontroller101 <= 64'd0;
		mem_ctrl_memorycontroller102 <= 64'd0;
		mem_ctrl_memorycontroller103 <= 64'd0;
		mem_ctrl_memorycontroller104 <= 64'd0;
		mem_ctrl_memorycontroller105 <= 64'd0;
		mem_ctrl_memorycontroller106 <= 64'd0;
		mem_ctrl_memorycontroller107 <= 64'd0;
		mem_ctrl_memorycontroller108 <= 64'd0;
		mem_ctrl_memorycontroller109 <= 64'd0;
		mem_ctrl_memorycontroller110 <= 64'd0;
		mem_ctrl_memorycontroller111 <= 64'd0;
		mem_ctrl_memorycontroller112 <= 64'd0;
		mem_ctrl_memorycontroller113 <= 64'd0;
		mem_ctrl_memorycontroller114 <= 64'd0;
		mem_ctrl_memorycontroller115 <= 64'd0;
		mem_ctrl_memorycontroller116 <= 64'd0;
		mem_ctrl_memorycontroller117 <= 64'd0;
		mem_ctrl_memorycontroller118 <= 64'd0;
		mem_ctrl_memorycontroller119 <= 64'd0;
		mem_ctrl_memorycontroller120 <= 64'd0;
		mem_ctrl_memorycontroller121 <= 64'd0;
		mem_ctrl_memorycontroller122 <= 64'd0;
		mem_ctrl_memorycontroller123 <= 64'd0;
		mem_ctrl_memorycontroller124 <= 64'd0;
		mem_ctrl_memorycontroller125 <= 64'd0;
		mem_ctrl_memorycontroller126 <= 64'd0;
		mem_ctrl_memorycontroller127 <= 64'd0;
		mem_ctrl_memorycontroller128 <= 64'd0;
		mem_ctrl_memorycontroller129 <= 64'd0;
		mem_ctrl_memorycontroller130 <= 64'd0;
		mem_ctrl_memorycontroller131 <= 64'd0;
		mem_ctrl_memorycontroller132 <= 64'd0;
		mem_ctrl_memorycontroller133 <= 64'd0;
		mem_ctrl_memorycontroller134 <= 64'd0;
		mem_ctrl_memorycontroller135 <= 64'd0;
		mem_ctrl_memorycontroller136 <= 64'd0;
		mem_ctrl_memorycontroller137 <= 64'd0;
		mem_ctrl_memorycontroller138 <= 64'd0;
		mem_ctrl_memorycontroller139 <= 64'd0;
		mem_ctrl_memorycontroller140 <= 64'd0;
		mem_ctrl_memorycontroller141 <= 64'd0;
		mem_ctrl_memorycontroller142 <= 64'd0;
		mem_ctrl_memorycontroller143 <= 64'd0;
		mem_ctrl_memorycontroller144 <= 64'd0;
		mem_ctrl_memorycontroller145 <= 64'd0;
		mem_ctrl_memorycontroller146 <= 64'd0;
		mem_ctrl_memorycontroller147 <= 64'd0;
		mem_ctrl_memorycontroller148 <= 64'd0;
		mem_ctrl_memorycontroller149 <= 64'd0;
		mem_ctrl_memorycontroller150 <= 64'd0;
		mem_ctrl_memorycontroller151 <= 64'd0;
		mem_ctrl_memorycontroller152 <= 64'd0;
		mem_ctrl_memorycontroller153 <= 64'd0;
		mem_ctrl_memorycontroller154 <= 64'd0;
		mem_ctrl_memorycontroller155 <= 64'd0;
		mem_ctrl_memorycontroller156 <= 64'd0;
		mem_ctrl_memorycontroller157 <= 64'd0;
		mem_ctrl_memorycontroller158 <= 64'd0;
		mem_ctrl_memorycontroller159 <= 64'd0;
		mem_ctrl_memorycontroller160 <= 64'd0;
		mem_ctrl_memorycontroller161 <= 64'd0;
		mem_ctrl_memorycontroller162 <= 64'd0;
		mem_ctrl_memorycontroller163 <= 64'd0;
		mem_ctrl_memorycontroller164 <= 64'd0;
		mem_ctrl_memorycontroller165 <= 64'd0;
		mem_ctrl_memorycontroller166 <= 64'd0;
		mem_ctrl_memorycontroller167 <= 64'd0;
		mem_ctrl_memorycontroller168 <= 64'd0;
		mem_ctrl_memorycontroller169 <= 64'd0;
		mem_ctrl_memorycontroller170 <= 64'd0;
		mem_ctrl_memorycontroller171 <= 64'd0;
		mem_ctrl_memorycontroller172 <= 64'd0;
		mem_ctrl_memorycontroller173 <= 64'd0;
		mem_ctrl_memorycontroller174 <= 64'd0;
		mem_ctrl_memorycontroller175 <= 64'd0;
		mem_ctrl_memorycontroller176 <= 64'd0;
		mem_ctrl_memorycontroller177 <= 64'd0;
		mem_ctrl_memorycontroller178 <= 64'd0;
		mem_ctrl_memorycontroller179 <= 64'd0;
		mem_ctrl_memorycontroller180 <= 64'd0;
		mem_ctrl_memorycontroller181 <= 64'd0;
		mem_ctrl_memorycontroller182 <= 64'd0;
		mem_ctrl_memorycontroller183 <= 64'd0;
		mem_ctrl_memorycontroller184 <= 64'd0;
		mem_ctrl_memorycontroller185 <= 64'd0;
		mem_ctrl_memorycontroller186 <= 64'd0;
		mem_ctrl_memorycontroller187 <= 64'd0;
		mem_ctrl_memorycontroller188 <= 64'd0;
		mem_ctrl_memorycontroller189 <= 64'd0;
		mem_ctrl_memorycontroller190 <= 64'd0;
		mem_ctrl_memorycontroller191 <= 64'd0;
		mem_ctrl_memorycontroller192 <= 64'd0;
		mem_ctrl_memorycontroller193 <= 64'd0;
		mem_ctrl_memorycontroller194 <= 64'd0;
		mem_ctrl_memorycontroller195 <= 64'd0;
		mem_ctrl_memorycontroller196 <= 64'd0;
		mem_ctrl_memorycontroller197 <= 64'd0;
		mem_ctrl_memorycontroller198 <= 64'd0;
		mem_ctrl_memorycontroller199 <= 64'd0;
		mem_ctrl_memorycontroller200 <= 64'd0;
		mem_ctrl_memorycontroller201 <= 64'd0;
		mem_ctrl_memorycontroller202 <= 64'd0;
		mem_ctrl_memorycontroller203 <= 64'd0;
		mem_ctrl_memorycontroller204 <= 64'd0;
		mem_ctrl_memorycontroller205 <= 64'd0;
		mem_ctrl_memorycontroller206 <= 64'd0;
		mem_ctrl_memorycontroller207 <= 64'd0;
		mem_ctrl_memorycontroller208 <= 64'd0;
		mem_ctrl_memorycontroller209 <= 64'd0;
		mem_ctrl_memorycontroller210 <= 64'd0;
		mem_ctrl_memorycontroller211 <= 64'd0;
		mem_ctrl_memorycontroller212 <= 64'd0;
		mem_ctrl_memorycontroller213 <= 64'd0;
		mem_ctrl_memorycontroller214 <= 64'd0;
		mem_ctrl_memorycontroller215 <= 64'd0;
		mem_ctrl_memorycontroller216 <= 64'd0;
		mem_ctrl_memorycontroller217 <= 64'd0;
		mem_ctrl_memorycontroller218 <= 64'd0;
		mem_ctrl_memorycontroller219 <= 64'd0;
		mem_ctrl_memorycontroller220 <= 64'd0;
		mem_ctrl_memorycontroller221 <= 64'd0;
		mem_ctrl_memorycontroller222 <= 64'd0;
		mem_ctrl_memorycontroller223 <= 64'd0;
		mem_ctrl_memorycontroller224 <= 64'd0;
		mem_ctrl_memorycontroller225 <= 64'd0;
		mem_ctrl_memorycontroller226 <= 64'd0;
		mem_ctrl_memorycontroller227 <= 64'd0;
		mem_ctrl_memorycontroller228 <= 64'd0;
		mem_ctrl_memorycontroller229 <= 64'd0;
		mem_ctrl_memorycontroller230 <= 64'd0;
		mem_ctrl_memorycontroller231 <= 64'd0;
		mem_ctrl_memorycontroller232 <= 64'd0;
		mem_ctrl_memorycontroller233 <= 64'd0;
		mem_ctrl_memorycontroller234 <= 64'd0;
		mem_ctrl_memorycontroller235 <= 64'd0;
		mem_ctrl_memorycontroller236 <= 64'd0;
		mem_ctrl_memorycontroller237 <= 64'd0;
		mem_ctrl_memorycontroller238 <= 64'd0;
		mem_ctrl_memorycontroller239 <= 64'd0;
		mem_ctrl_memorycontroller240 <= 64'd0;
		mem_ctrl_memorycontroller241 <= 64'd0;
		mem_ctrl_memorycontroller242 <= 64'd0;
		mem_ctrl_memorycontroller243 <= 64'd0;
		mem_ctrl_memorycontroller244 <= 64'd0;
		mem_ctrl_memorycontroller245 <= 64'd0;
		mem_ctrl_memorycontroller246 <= 64'd0;
		mem_ctrl_memorycontroller247 <= 64'd0;
		mem_ctrl_memorycontroller248 <= 64'd0;
		mem_ctrl_memorycontroller249 <= 64'd0;
		mem_ctrl_memorycontroller250 <= 64'd0;
		mem_ctrl_memorycontroller251 <= 64'd0;
		mem_ctrl_memorycontroller252 <= 64'd0;
		mem_ctrl_memorycontroller253 <= 64'd0;
		mem_ctrl_memorycontroller254 <= 64'd0;
		mem_ctrl_memorycontroller255 <= 64'd0;
		mem_ctrl_memorycontroller256 <= 64'd0;
		mem_ctrl_memorycontroller257 <= 64'd0;
		mem_ctrl_memorycontroller258 <= 64'd0;
		mem_ctrl_memorycontroller259 <= 64'd0;
		mem_ctrl_memorycontroller260 <= 64'd0;
		mem_ctrl_memorycontroller261 <= 64'd0;
		mem_ctrl_memorycontroller262 <= 64'd0;
		mem_ctrl_memorycontroller263 <= 64'd0;
		mem_ctrl_memorycontroller264 <= 64'd0;
		mem_ctrl_memorycontroller265 <= 64'd0;
		mem_ctrl_memorycontroller266 <= 64'd0;
		mem_ctrl_memorycontroller267 <= 64'd0;
		mem_ctrl_memorycontroller268 <= 64'd0;
		mem_ctrl_memorycontroller269 <= 64'd0;
		mem_ctrl_memorycontroller270 <= 64'd0;
		mem_ctrl_memorycontroller271 <= 64'd0;
		mem_ctrl_memorycontroller272 <= 64'd0;
		mem_ctrl_memorycontroller273 <= 64'd0;
		mem_ctrl_memorycontroller274 <= 64'd0;
		mem_ctrl_memorycontroller275 <= 64'd0;
		mem_ctrl_memorycontroller276 <= 64'd0;
		mem_ctrl_memorycontroller277 <= 64'd0;
		mem_ctrl_memorycontroller278 <= 64'd0;
		mem_ctrl_memorycontroller279 <= 64'd0;
		mem_ctrl_memorycontroller280 <= 64'd0;
		mem_ctrl_memorycontroller281 <= 64'd0;
		mem_ctrl_memorycontroller282 <= 64'd0;
		mem_ctrl_memorycontroller283 <= 64'd0;
		mem_ctrl_memorycontroller284 <= 64'd0;
		mem_ctrl_memorycontroller285 <= 64'd0;
		mem_ctrl_memorycontroller286 <= 64'd0;
		mem_ctrl_memorycontroller287 <= 64'd0;
		mem_ctrl_memorycontroller288 <= 64'd0;
		mem_ctrl_memorycontroller289 <= 64'd0;
		mem_ctrl_memorycontroller290 <= 64'd0;
		mem_ctrl_memorycontroller291 <= 64'd0;
		mem_ctrl_memorycontroller292 <= 64'd0;
		mem_ctrl_memorycontroller293 <= 64'd0;
		mem_ctrl_memorycontroller294 <= 64'd0;
		mem_ctrl_memorycontroller295 <= 64'd0;
		mem_ctrl_memorycontroller296 <= 64'd0;
		mem_ctrl_memorycontroller297 <= 64'd0;
		mem_ctrl_memorycontroller298 <= 64'd0;
		mem_ctrl_memorycontroller299 <= 64'd0;
		mem_ctrl_memorycontroller300 <= 64'd0;
		mem_ctrl_memorycontroller301 <= 64'd0;
		mem_ctrl_memorycontroller302 <= 64'd0;
		mem_ctrl_memorycontroller303 <= 64'd0;
		mem_ctrl_memorycontroller304 <= 64'd0;
		mem_ctrl_memorycontroller305 <= 64'd0;
		mem_ctrl_memorycontroller306 <= 64'd0;
		mem_ctrl_memorycontroller307 <= 64'd0;
		mem_ctrl_memorycontroller308 <= 64'd0;
		mem_ctrl_memorycontroller309 <= 64'd0;
		mem_ctrl_memorycontroller310 <= 64'd0;
		mem_ctrl_memorycontroller311 <= 64'd0;
		mem_ctrl_memorycontroller312 <= 64'd0;
		mem_ctrl_memorycontroller313 <= 64'd0;
		mem_ctrl_memorycontroller314 <= 64'd0;
		mem_ctrl_memorycontroller315 <= 64'd0;
		mem_ctrl_memorycontroller316 <= 64'd0;
		mem_ctrl_memorycontroller317 <= 64'd0;
		mem_ctrl_memorycontroller318 <= 64'd0;
		mem_ctrl_memorycontroller319 <= 64'd0;
		mem_ctrl_memorycontroller320 <= 64'd0;
		mem_ctrl_memorycontroller321 <= 64'd0;
		mem_ctrl_memorycontroller322 <= 64'd0;
		mem_ctrl_memorycontroller323 <= 64'd0;
		mem_ctrl_memorycontroller324 <= 64'd0;
		mem_ctrl_memorycontroller325 <= 64'd0;
		mem_ctrl_memorycontroller326 <= 64'd0;
		mem_ctrl_memorycontroller327 <= 64'd0;
		mem_ctrl_memorycontroller328 <= 64'd0;
		mem_ctrl_memorycontroller329 <= 64'd0;
		mem_ctrl_memorycontroller330 <= 64'd0;
		mem_ctrl_memorycontroller331 <= 64'd0;
		mem_ctrl_memorycontroller332 <= 64'd0;
		mem_ctrl_memorycontroller333 <= 64'd0;
		mem_ctrl_memorycontroller334 <= 64'd0;
		mem_ctrl_memorycontroller335 <= 64'd0;
		mem_ctrl_memorycontroller336 <= 64'd0;
		mem_ctrl_memorycontroller337 <= 64'd0;
		mem_ctrl_memorycontroller338 <= 64'd0;
		mem_ctrl_memorycontroller339 <= 64'd0;
		mem_ctrl_memorycontroller340 <= 64'd0;
		mem_ctrl_memorycontroller341 <= 64'd0;
		mem_ctrl_memorycontroller342 <= 64'd0;
		mem_ctrl_memorycontroller343 <= 64'd0;
		mem_ctrl_memorycontroller344 <= 64'd0;
		mem_ctrl_memorycontroller345 <= 64'd0;
		mem_ctrl_memorycontroller346 <= 64'd0;
		mem_ctrl_memorycontroller347 <= 64'd0;
		mem_ctrl_memorycontroller348 <= 64'd0;
		mem_ctrl_memorycontroller349 <= 64'd0;
		mem_ctrl_memorycontroller350 <= 64'd0;
		mem_ctrl_memorycontroller351 <= 64'd0;
		mem_ctrl_memorycontroller352 <= 64'd0;
		mem_ctrl_memorycontroller353 <= 64'd0;
		mem_ctrl_memorycontroller354 <= 64'd0;
		mem_ctrl_memorycontroller355 <= 64'd0;
		mem_ctrl_memorycontroller356 <= 64'd0;
		mem_ctrl_memorycontroller357 <= 64'd0;
		mem_ctrl_memorycontroller358 <= 64'd0;
		mem_ctrl_memorycontroller359 <= 64'd0;
		mem_ctrl_memorycontroller360 <= 64'd0;
		mem_ctrl_memorycontroller361 <= 64'd0;
		mem_ctrl_memorycontroller362 <= 64'd0;
		mem_ctrl_memorycontroller363 <= 64'd0;
		mem_ctrl_memorycontroller364 <= 64'd0;
		mem_ctrl_memorycontroller365 <= 64'd0;
		mem_ctrl_memorycontroller366 <= 64'd0;
		mem_ctrl_memorycontroller367 <= 64'd0;
		mem_ctrl_memorycontroller368 <= 64'd0;
		mem_ctrl_memorycontroller369 <= 64'd0;
		mem_ctrl_memorycontroller370 <= 64'd0;
		mem_ctrl_memorycontroller371 <= 64'd0;
		mem_ctrl_memorycontroller372 <= 64'd0;
		mem_ctrl_memorycontroller373 <= 64'd0;
		mem_ctrl_memorycontroller374 <= 64'd0;
		mem_ctrl_memorycontroller375 <= 64'd0;
		mem_ctrl_memorycontroller376 <= 64'd0;
		mem_ctrl_memorycontroller377 <= 64'd0;
		mem_ctrl_memorycontroller378 <= 64'd0;
		mem_ctrl_memorycontroller379 <= 64'd0;
		mem_ctrl_memorycontroller380 <= 64'd0;
		mem_ctrl_memorycontroller381 <= 64'd0;
		mem_ctrl_memorycontroller382 <= 64'd0;
		mem_ctrl_memorycontroller383 <= 64'd0;
		mem_ctrl_memorycontroller384 <= 64'd0;
		mem_ctrl_memorycontroller385 <= 64'd0;
		mem_ctrl_memorycontroller386 <= 64'd0;
		mem_ctrl_memorycontroller387 <= 64'd0;
		mem_ctrl_memorycontroller388 <= 64'd0;
		mem_ctrl_memorycontroller389 <= 64'd0;
		mem_ctrl_memorycontroller390 <= 64'd0;
		mem_ctrl_memorycontroller391 <= 64'd0;
		mem_ctrl_memorycontroller392 <= 64'd0;
		mem_ctrl_memorycontroller393 <= 64'd0;
		mem_ctrl_memorycontroller394 <= 64'd0;
		mem_ctrl_memorycontroller395 <= 64'd0;
		mem_ctrl_memorycontroller396 <= 64'd0;
		mem_ctrl_memorycontroller397 <= 64'd0;
		mem_ctrl_memorycontroller398 <= 64'd0;
		mem_ctrl_memorycontroller399 <= 64'd0;
		mem_ctrl_memorycontroller400 <= 64'd0;
		mem_ctrl_memorycontroller401 <= 64'd0;
		mem_ctrl_memorycontroller402 <= 64'd0;
		mem_ctrl_memorycontroller403 <= 64'd0;
		mem_ctrl_memorycontroller404 <= 64'd0;
		mem_ctrl_memorycontroller405 <= 64'd0;
		mem_ctrl_memorycontroller406 <= 64'd0;
		mem_ctrl_memorycontroller407 <= 64'd0;
		mem_ctrl_memorycontroller408 <= 64'd0;
		mem_ctrl_memorycontroller409 <= 64'd0;
		mem_ctrl_memorycontroller410 <= 64'd0;
		mem_ctrl_memorycontroller411 <= 64'd0;
		mem_ctrl_memorycontroller412 <= 64'd0;
		mem_ctrl_memorycontroller413 <= 64'd0;
		mem_ctrl_memorycontroller414 <= 64'd0;
		mem_ctrl_memorycontroller415 <= 64'd0;
		mem_ctrl_memorycontroller416 <= 64'd0;
		mem_ctrl_memorycontroller417 <= 64'd0;
		mem_ctrl_memorycontroller418 <= 64'd0;
		mem_ctrl_memorycontroller419 <= 64'd0;
		mem_ctrl_memorycontroller420 <= 64'd0;
		mem_ctrl_memorycontroller421 <= 64'd0;
		mem_ctrl_memorycontroller422 <= 64'd0;
		mem_ctrl_memorycontroller423 <= 64'd0;
		mem_ctrl_memorycontroller424 <= 64'd0;
		mem_ctrl_memorycontroller425 <= 64'd0;
		mem_ctrl_memorycontroller426 <= 64'd0;
		mem_ctrl_memorycontroller427 <= 64'd0;
		mem_ctrl_memorycontroller428 <= 64'd0;
		mem_ctrl_memorycontroller429 <= 64'd0;
		mem_ctrl_memorycontroller430 <= 64'd0;
		mem_ctrl_memorycontroller431 <= 64'd0;
		mem_ctrl_memorycontroller432 <= 64'd0;
		mem_ctrl_memorycontroller433 <= 64'd0;
		mem_ctrl_memorycontroller434 <= 64'd0;
		mem_ctrl_memorycontroller435 <= 64'd0;
		mem_ctrl_memorycontroller436 <= 64'd0;
		mem_ctrl_memorycontroller437 <= 64'd0;
		mem_ctrl_memorycontroller438 <= 64'd0;
		mem_ctrl_memorycontroller439 <= 64'd0;
		mem_ctrl_memorycontroller440 <= 64'd0;
		mem_ctrl_memorycontroller441 <= 64'd0;
		mem_ctrl_memorycontroller442 <= 64'd0;
		mem_ctrl_memorycontroller443 <= 64'd0;
		mem_ctrl_memorycontroller444 <= 64'd0;
		mem_ctrl_memorycontroller445 <= 64'd0;
		mem_ctrl_memorycontroller446 <= 64'd0;
		mem_ctrl_memorycontroller447 <= 64'd0;
		mem_ctrl_memorycontroller448 <= 64'd0;
		mem_ctrl_memorycontroller449 <= 64'd0;
		mem_ctrl_memorycontroller450 <= 64'd0;
		mem_ctrl_memorycontroller451 <= 64'd0;
		mem_ctrl_memorycontroller452 <= 64'd0;
		mem_ctrl_memorycontroller453 <= 64'd0;
		mem_ctrl_memorycontroller454 <= 64'd0;
		mem_ctrl_memorycontroller455 <= 64'd0;
		mem_ctrl_memorycontroller456 <= 64'd0;
		mem_ctrl_memorycontroller457 <= 64'd0;
		mem_ctrl_memorycontroller458 <= 64'd0;
		mem_ctrl_memorycontroller459 <= 64'd0;
		mem_ctrl_memorycontroller460 <= 64'd0;
		mem_ctrl_memorycontroller461 <= 64'd0;
		mem_ctrl_memorycontroller462 <= 64'd0;
		mem_ctrl_memorycontroller463 <= 64'd0;
		mem_ctrl_memorycontroller464 <= 64'd0;
		mem_ctrl_memorycontroller465 <= 64'd0;
		mem_ctrl_memorycontroller466 <= 64'd0;
		mem_ctrl_memorycontroller467 <= 64'd0;
		mem_ctrl_memorycontroller468 <= 64'd0;
		mem_ctrl_memorycontroller469 <= 64'd0;
		mem_ctrl_memorycontroller470 <= 64'd0;
		mem_ctrl_memorycontroller471 <= 64'd0;
		mem_ctrl_memorycontroller472 <= 64'd0;
		mem_ctrl_memorycontroller473 <= 64'd0;
		mem_ctrl_memorycontroller474 <= 64'd0;
		mem_ctrl_memorycontroller475 <= 64'd0;
		mem_ctrl_memorycontroller476 <= 64'd0;
		mem_ctrl_memorycontroller477 <= 64'd0;
		mem_ctrl_memorycontroller478 <= 64'd0;
		mem_ctrl_memorycontroller479 <= 64'd0;
		mem_ctrl_memorycontroller480 <= 64'd0;
		mem_ctrl_memorycontroller481 <= 64'd0;
		mem_ctrl_memorycontroller482 <= 64'd0;
		mem_ctrl_memorycontroller483 <= 64'd0;
		mem_ctrl_memorycontroller484 <= 64'd0;
		mem_ctrl_memorycontroller485 <= 64'd0;
		mem_ctrl_memorycontroller486 <= 64'd0;
		mem_ctrl_memorycontroller487 <= 64'd0;
		mem_ctrl_memorycontroller488 <= 64'd0;
		mem_ctrl_memorycontroller489 <= 64'd0;
		mem_ctrl_memorycontroller490 <= 64'd0;
		mem_ctrl_memorycontroller491 <= 64'd0;
		mem_ctrl_memorycontroller492 <= 64'd0;
		mem_ctrl_memorycontroller493 <= 64'd0;
		mem_ctrl_memorycontroller494 <= 64'd0;
		mem_ctrl_memorycontroller495 <= 64'd0;
		mem_ctrl_memorycontroller496 <= 64'd0;
		mem_ctrl_memorycontroller497 <= 64'd0;
		mem_ctrl_memorycontroller498 <= 64'd0;
		mem_ctrl_memorycontroller499 <= 64'd0;
		mem_ctrl_memorycontroller500 <= 64'd0;
		mem_ctrl_memorycontroller501 <= 64'd0;
		mem_ctrl_memorycontroller502 <= 64'd0;
		mem_ctrl_memorycontroller503 <= 64'd0;
		mem_ctrl_memorycontroller504 <= 64'd0;
		mem_ctrl_memorycontroller505 <= 64'd0;
		mem_ctrl_memorycontroller506 <= 64'd0;
		mem_ctrl_memorycontroller507 <= 64'd0;
		mem_ctrl_memorycontroller508 <= 64'd0;
		mem_ctrl_memorycontroller509 <= 64'd0;
		mem_ctrl_memorycontroller510 <= 64'd0;
		mem_ctrl_memorycontroller511 <= 64'd0;
		mem_ctrl_memorycontroller512 <= 64'd0;
		mem_ctrl_memorycontroller513 <= 64'd0;
		mem_ctrl_memorycontroller514 <= 64'd0;
		mem_ctrl_memorycontroller515 <= 64'd0;
		mem_ctrl_memorycontroller516 <= 64'd0;
		mem_ctrl_memorycontroller517 <= 64'd0;
		mem_ctrl_memorycontroller518 <= 64'd0;
		mem_ctrl_memorycontroller519 <= 64'd0;
		mem_ctrl_memorycontroller520 <= 64'd0;
		mem_ctrl_memorycontroller521 <= 64'd0;
		mem_ctrl_memorycontroller522 <= 64'd0;
		mem_ctrl_memorycontroller523 <= 64'd0;
		mem_ctrl_memorycontroller524 <= 64'd0;
		mem_ctrl_memorycontroller525 <= 64'd0;
		mem_ctrl_memorycontroller526 <= 64'd0;
		mem_ctrl_memorycontroller527 <= 64'd0;
		mem_ctrl_memorycontroller528 <= 64'd0;
		mem_ctrl_memorycontroller529 <= 64'd0;
		mem_ctrl_memorycontroller530 <= 64'd0;
		mem_ctrl_memorycontroller531 <= 64'd0;
		mem_ctrl_memorycontroller532 <= 64'd0;
		mem_ctrl_memorycontroller533 <= 64'd0;
		mem_ctrl_memorycontroller534 <= 64'd0;
		mem_ctrl_memorycontroller535 <= 64'd0;
		mem_ctrl_memorycontroller536 <= 64'd0;
		mem_ctrl_memorycontroller537 <= 64'd0;
		mem_ctrl_memorycontroller538 <= 64'd0;
		mem_ctrl_memorycontroller539 <= 64'd0;
		mem_ctrl_memorycontroller540 <= 64'd0;
		mem_ctrl_memorycontroller541 <= 64'd0;
		mem_ctrl_memorycontroller542 <= 64'd0;
		mem_ctrl_memorycontroller543 <= 64'd0;
		mem_ctrl_memorycontroller544 <= 64'd0;
		mem_ctrl_memorycontroller545 <= 64'd0;
		mem_ctrl_memorycontroller546 <= 64'd0;
		mem_ctrl_memorycontroller547 <= 64'd0;
		mem_ctrl_memorycontroller548 <= 64'd0;
		mem_ctrl_memorycontroller549 <= 64'd0;
		mem_ctrl_memorycontroller550 <= 64'd0;
		mem_ctrl_memorycontroller551 <= 64'd0;
		mem_ctrl_memorycontroller552 <= 64'd0;
		mem_ctrl_memorycontroller553 <= 64'd0;
		mem_ctrl_memorycontroller554 <= 64'd0;
		mem_ctrl_memorycontroller555 <= 64'd0;
		mem_ctrl_memorycontroller556 <= 64'd0;
		mem_ctrl_memorycontroller557 <= 64'd0;
		mem_ctrl_memorycontroller558 <= 64'd0;
		mem_ctrl_memorycontroller559 <= 64'd0;
		mem_ctrl_memorycontroller560 <= 64'd0;
		mem_ctrl_memorycontroller561 <= 64'd0;
		mem_ctrl_memorycontroller562 <= 64'd0;
		mem_ctrl_memorycontroller563 <= 64'd0;
		mem_ctrl_memorycontroller564 <= 64'd0;
		mem_ctrl_memorycontroller565 <= 64'd0;
		mem_ctrl_memorycontroller566 <= 64'd0;
		mem_ctrl_memorycontroller567 <= 64'd0;
		mem_ctrl_memorycontroller568 <= 64'd0;
		mem_ctrl_memorycontroller569 <= 64'd0;
		mem_ctrl_memorycontroller570 <= 64'd0;
		mem_ctrl_memorycontroller571 <= 64'd0;
		mem_ctrl_memorycontroller572 <= 64'd0;
		mem_ctrl_memorycontroller573 <= 64'd0;
		mem_ctrl_memorycontroller574 <= 64'd0;
		mem_ctrl_memorycontroller575 <= 64'd0;
		mem_ctrl_memorycontroller576 <= 64'd0;
		mem_ctrl_memorycontroller577 <= 64'd0;
		mem_ctrl_memorycontroller578 <= 64'd0;
		mem_ctrl_memorycontroller579 <= 64'd0;
		mem_ctrl_memorycontroller580 <= 64'd0;
		mem_ctrl_memorycontroller581 <= 64'd0;
		mem_ctrl_memorycontroller582 <= 64'd0;
		mem_ctrl_memorycontroller583 <= 64'd0;
		mem_ctrl_memorycontroller584 <= 64'd0;
		mem_ctrl_memorycontroller585 <= 64'd0;
		mem_ctrl_memorycontroller586 <= 64'd0;
		mem_ctrl_memorycontroller587 <= 64'd0;
		mem_ctrl_memorycontroller588 <= 64'd0;
		mem_ctrl_memorycontroller589 <= 64'd0;
		mem_ctrl_memorycontroller590 <= 64'd0;
		mem_ctrl_memorycontroller591 <= 64'd0;
		mem_ctrl_memorycontroller592 <= 64'd0;
		mem_ctrl_memorycontroller593 <= 64'd0;
		mem_ctrl_memorycontroller594 <= 64'd0;
		mem_ctrl_memorycontroller595 <= 64'd0;
		mem_ctrl_memorycontroller596 <= 64'd0;
		mem_ctrl_memorycontroller597 <= 64'd0;
		mem_ctrl_memorycontroller598 <= 64'd0;
		mem_ctrl_memorycontroller599 <= 64'd0;
		mem_ctrl_memorycontroller600 <= 64'd0;
		mem_ctrl_memorycontroller601 <= 64'd0;
		mem_ctrl_memorycontroller602 <= 64'd0;
		mem_ctrl_memorycontroller603 <= 64'd0;
		mem_ctrl_memorycontroller604 <= 64'd0;
		mem_ctrl_memorycontroller605 <= 64'd0;
		mem_ctrl_memorycontroller606 <= 64'd0;
		mem_ctrl_memorycontroller607 <= 64'd0;
		mem_ctrl_memorycontroller608 <= 64'd0;
		mem_ctrl_memorycontroller609 <= 64'd0;
		mem_ctrl_memorycontroller610 <= 64'd0;
		mem_ctrl_memorycontroller611 <= 64'd0;
		mem_ctrl_memorycontroller612 <= 64'd0;
		mem_ctrl_memorycontroller613 <= 64'd0;
		mem_ctrl_memorycontroller614 <= 64'd0;
		mem_ctrl_memorycontroller615 <= 64'd0;
		mem_ctrl_memorycontroller616 <= 64'd0;
		mem_ctrl_memorycontroller617 <= 64'd0;
		mem_ctrl_memorycontroller618 <= 64'd0;
		mem_ctrl_memorycontroller619 <= 64'd0;
		mem_ctrl_memorycontroller620 <= 64'd0;
		mem_ctrl_memorycontroller621 <= 64'd0;
		mem_ctrl_memorycontroller622 <= 64'd0;
		mem_ctrl_memorycontroller623 <= 64'd0;
		mem_ctrl_memorycontroller624 <= 64'd0;
		mem_ctrl_memorycontroller625 <= 64'd0;
		mem_ctrl_memorycontroller626 <= 64'd0;
		mem_ctrl_memorycontroller627 <= 64'd0;
		mem_ctrl_memorycontroller628 <= 64'd0;
		mem_ctrl_memorycontroller629 <= 64'd0;
		mem_ctrl_memorycontroller630 <= 64'd0;
		mem_ctrl_memorycontroller631 <= 64'd0;
		mem_ctrl_memorycontroller632 <= 64'd0;
		mem_ctrl_memorycontroller633 <= 64'd0;
		mem_ctrl_memorycontroller634 <= 64'd0;
		mem_ctrl_memorycontroller635 <= 64'd0;
		mem_ctrl_memorycontroller636 <= 64'd0;
		mem_ctrl_memorycontroller637 <= 64'd0;
		mem_ctrl_memorycontroller638 <= 64'd0;
		mem_ctrl_memorycontroller639 <= 64'd0;
		mem_ctrl_memorycontroller640 <= 64'd0;
		mem_ctrl_memorycontroller641 <= 64'd0;
		mem_ctrl_memorycontroller642 <= 64'd0;
		mem_ctrl_memorycontroller643 <= 64'd0;
		mem_ctrl_memorycontroller644 <= 64'd0;
		mem_ctrl_memorycontroller645 <= 64'd0;
		mem_ctrl_memorycontroller646 <= 64'd0;
		mem_ctrl_memorycontroller647 <= 64'd0;
		mem_ctrl_memorycontroller648 <= 64'd0;
		mem_ctrl_memorycontroller649 <= 64'd0;
		mem_ctrl_memorycontroller650 <= 64'd0;
		mem_ctrl_memorycontroller651 <= 64'd0;
		mem_ctrl_memorycontroller652 <= 64'd0;
		mem_ctrl_memorycontroller653 <= 64'd0;
		mem_ctrl_memorycontroller654 <= 64'd0;
		mem_ctrl_memorycontroller655 <= 64'd0;
		mem_ctrl_memorycontroller656 <= 64'd0;
		mem_ctrl_memorycontroller657 <= 64'd0;
		mem_ctrl_memorycontroller658 <= 64'd0;
		mem_ctrl_memorycontroller659 <= 64'd0;
		mem_ctrl_memorycontroller660 <= 64'd0;
		mem_ctrl_memorycontroller661 <= 64'd0;
		mem_ctrl_memorycontroller662 <= 64'd0;
		mem_ctrl_memorycontroller663 <= 64'd0;
		mem_ctrl_memorycontroller664 <= 64'd0;
		mem_ctrl_memorycontroller665 <= 64'd0;
		mem_ctrl_memorycontroller666 <= 64'd0;
		mem_ctrl_memorycontroller667 <= 64'd0;
		mem_ctrl_memorycontroller668 <= 64'd0;
		mem_ctrl_memorycontroller669 <= 64'd0;
		mem_ctrl_memorycontroller670 <= 64'd0;
		mem_ctrl_memorycontroller671 <= 64'd0;
		mem_ctrl_memorycontroller672 <= 64'd0;
		mem_ctrl_memorycontroller673 <= 64'd0;
		mem_ctrl_memorycontroller674 <= 64'd0;
		mem_ctrl_memorycontroller675 <= 64'd0;
		mem_ctrl_memorycontroller676 <= 64'd0;
		mem_ctrl_memorycontroller677 <= 64'd0;
		mem_ctrl_memorycontroller678 <= 64'd0;
		mem_ctrl_memorycontroller679 <= 64'd0;
		mem_ctrl_memorycontroller680 <= 64'd0;
		mem_ctrl_memorycontroller681 <= 64'd0;
		mem_ctrl_memorycontroller682 <= 64'd0;
		mem_ctrl_memorycontroller683 <= 64'd0;
		mem_ctrl_memorycontroller684 <= 64'd0;
		mem_ctrl_memorycontroller685 <= 64'd0;
		mem_ctrl_memorycontroller686 <= 64'd0;
		mem_ctrl_memorycontroller687 <= 64'd0;
		mem_ctrl_memorycontroller688 <= 64'd0;
		mem_ctrl_memorycontroller689 <= 64'd0;
		mem_ctrl_memorycontroller690 <= 64'd0;
		mem_ctrl_memorycontroller691 <= 64'd0;
		mem_ctrl_memorycontroller692 <= 64'd0;
		mem_ctrl_memorycontroller693 <= 64'd0;
		mem_ctrl_memorycontroller694 <= 64'd0;
		mem_ctrl_memorycontroller695 <= 64'd0;
		mem_ctrl_memorycontroller696 <= 64'd0;
		mem_ctrl_memorycontroller697 <= 64'd0;
		mem_ctrl_memorycontroller698 <= 64'd0;
		mem_ctrl_memorycontroller699 <= 64'd0;
		mem_ctrl_memorycontroller700 <= 64'd0;
		mem_ctrl_memorycontroller701 <= 64'd0;
		mem_ctrl_memorycontroller702 <= 64'd0;
		mem_ctrl_memorycontroller703 <= 64'd0;
		mem_ctrl_memorycontroller704 <= 64'd0;
		mem_ctrl_memorycontroller705 <= 64'd0;
		mem_ctrl_memorycontroller706 <= 64'd0;
		mem_ctrl_memorycontroller707 <= 64'd0;
		mem_ctrl_memorycontroller708 <= 64'd0;
		mem_ctrl_memorycontroller709 <= 64'd0;
		mem_ctrl_memorycontroller710 <= 64'd0;
		mem_ctrl_memorycontroller711 <= 64'd0;
		mem_ctrl_memorycontroller712 <= 64'd0;
		mem_ctrl_memorycontroller713 <= 64'd0;
		mem_ctrl_memorycontroller714 <= 64'd0;
		mem_ctrl_memorycontroller715 <= 64'd0;
		mem_ctrl_memorycontroller716 <= 64'd0;
		mem_ctrl_memorycontroller717 <= 64'd0;
		mem_ctrl_memorycontroller718 <= 64'd0;
		mem_ctrl_memorycontroller719 <= 64'd0;
		mem_ctrl_memorycontroller720 <= 64'd0;
		mem_ctrl_memorycontroller721 <= 64'd0;
		mem_ctrl_memorycontroller722 <= 64'd0;
		mem_ctrl_memorycontroller723 <= 64'd0;
		mem_ctrl_memorycontroller724 <= 64'd0;
		mem_ctrl_memorycontroller725 <= 64'd0;
		mem_ctrl_memorycontroller726 <= 64'd0;
		mem_ctrl_memorycontroller727 <= 64'd0;
		mem_ctrl_memorycontroller728 <= 64'd0;
		mem_ctrl_memorycontroller729 <= 64'd0;
		mem_ctrl_memorycontroller730 <= 64'd0;
		mem_ctrl_memorycontroller731 <= 64'd0;
		mem_ctrl_memorycontroller732 <= 64'd0;
		mem_ctrl_memorycontroller733 <= 64'd0;
		mem_ctrl_memorycontroller734 <= 64'd0;
		mem_ctrl_memorycontroller735 <= 64'd0;
		mem_ctrl_memorycontroller736 <= 64'd0;
		mem_ctrl_memorycontroller737 <= 64'd0;
		mem_ctrl_memorycontroller738 <= 64'd0;
		mem_ctrl_memorycontroller739 <= 64'd0;
		mem_ctrl_memorycontroller740 <= 64'd0;
		mem_ctrl_memorycontroller741 <= 64'd0;
		mem_ctrl_memorycontroller742 <= 64'd0;
		mem_ctrl_memorycontroller743 <= 64'd0;
		mem_ctrl_memorycontroller744 <= 64'd0;
		mem_ctrl_memorycontroller745 <= 64'd0;
		mem_ctrl_memorycontroller746 <= 64'd0;
		mem_ctrl_memorycontroller747 <= 64'd0;
		mem_ctrl_memorycontroller748 <= 64'd0;
		mem_ctrl_memorycontroller749 <= 64'd0;
		mem_ctrl_memorycontroller750 <= 64'd0;
		mem_ctrl_memorycontroller751 <= 64'd0;
		mem_ctrl_memorycontroller752 <= 64'd0;
		mem_ctrl_memorycontroller753 <= 64'd0;
		mem_ctrl_memorycontroller754 <= 64'd0;
		mem_ctrl_memorycontroller755 <= 64'd0;
		mem_ctrl_memorycontroller756 <= 64'd0;
		mem_ctrl_memorycontroller757 <= 64'd0;
		mem_ctrl_memorycontroller758 <= 64'd0;
		mem_ctrl_memorycontroller759 <= 64'd0;
		mem_ctrl_memorycontroller760 <= 64'd0;
		mem_ctrl_memorycontroller761 <= 64'd0;
		mem_ctrl_memorycontroller762 <= 64'd0;
		mem_ctrl_memorycontroller763 <= 64'd0;
		mem_ctrl_memorycontroller764 <= 64'd0;
		mem_ctrl_memorycontroller765 <= 64'd0;
		mem_ctrl_memorycontroller766 <= 64'd0;
		mem_ctrl_memorycontroller767 <= 64'd0;
		mem_ctrl_memorycontroller768 <= 64'd0;
		mem_ctrl_memorycontroller769 <= 64'd0;
		mem_ctrl_memorycontroller770 <= 64'd0;
		mem_ctrl_memorycontroller771 <= 64'd0;
		mem_ctrl_memorycontroller772 <= 64'd0;
		mem_ctrl_memorycontroller773 <= 64'd0;
		mem_ctrl_memorycontroller774 <= 64'd0;
		mem_ctrl_memorycontroller775 <= 64'd0;
		mem_ctrl_memorycontroller776 <= 64'd0;
		mem_ctrl_memorycontroller777 <= 64'd0;
		mem_ctrl_memorycontroller778 <= 64'd0;
		mem_ctrl_memorycontroller779 <= 64'd0;
		mem_ctrl_memorycontroller780 <= 64'd0;
		mem_ctrl_memorycontroller781 <= 64'd0;
		mem_ctrl_memorycontroller782 <= 64'd0;
		mem_ctrl_memorycontroller783 <= 64'd0;
		mem_ctrl_memorycontroller784 <= 64'd0;
		mem_ctrl_memorycontroller785 <= 64'd0;
		mem_ctrl_memorycontroller786 <= 64'd0;
		mem_ctrl_memorycontroller787 <= 64'd0;
		mem_ctrl_memorycontroller788 <= 64'd0;
		mem_ctrl_memorycontroller789 <= 64'd0;
		mem_ctrl_memorycontroller790 <= 64'd0;
		mem_ctrl_memorycontroller791 <= 64'd0;
		mem_ctrl_memorycontroller792 <= 64'd0;
		mem_ctrl_memorycontroller793 <= 64'd0;
		mem_ctrl_memorycontroller794 <= 64'd0;
		mem_ctrl_memorycontroller795 <= 64'd0;
		mem_ctrl_memorycontroller796 <= 64'd0;
		mem_ctrl_memorycontroller797 <= 64'd0;
		mem_ctrl_memorycontroller798 <= 64'd0;
		mem_ctrl_memorycontroller799 <= 64'd0;
		mem_ctrl_memorycontroller800 <= 64'd0;
		mem_ctrl_memorycontroller801 <= 64'd0;
		mem_ctrl_memorycontroller802 <= 64'd0;
		mem_ctrl_memorycontroller803 <= 64'd0;
		mem_ctrl_memorycontroller804 <= 64'd0;
		mem_ctrl_memorycontroller805 <= 64'd0;
		mem_ctrl_memorycontroller806 <= 64'd0;
		mem_ctrl_memorycontroller807 <= 64'd0;
		mem_ctrl_memorycontroller808 <= 64'd0;
		mem_ctrl_memorycontroller809 <= 64'd0;
		mem_ctrl_memorycontroller810 <= 64'd0;
		mem_ctrl_memorycontroller811 <= 64'd0;
		mem_ctrl_memorycontroller812 <= 64'd0;
		mem_ctrl_memorycontroller813 <= 64'd0;
		mem_ctrl_memorycontroller814 <= 64'd0;
		mem_ctrl_memorycontroller815 <= 64'd0;
		mem_ctrl_memorycontroller816 <= 64'd0;
		mem_ctrl_memorycontroller817 <= 64'd0;
		mem_ctrl_memorycontroller818 <= 64'd0;
		mem_ctrl_memorycontroller819 <= 64'd0;
		mem_ctrl_memorycontroller820 <= 64'd0;
		mem_ctrl_memorycontroller821 <= 64'd0;
		mem_ctrl_memorycontroller822 <= 64'd0;
		mem_ctrl_memorycontroller823 <= 64'd0;
		mem_ctrl_memorycontroller824 <= 64'd0;
		mem_ctrl_memorycontroller825 <= 64'd0;
		mem_ctrl_memorycontroller826 <= 64'd0;
		mem_ctrl_memorycontroller827 <= 64'd0;
		mem_ctrl_memorycontroller828 <= 64'd0;
		mem_ctrl_memorycontroller829 <= 64'd0;
		mem_ctrl_memorycontroller830 <= 64'd0;
		mem_ctrl_memorycontroller831 <= 64'd0;
		mem_ctrl_memorycontroller832 <= 64'd0;
		mem_ctrl_memorycontroller833 <= 64'd0;
		mem_ctrl_memorycontroller834 <= 64'd0;
		mem_ctrl_memorycontroller835 <= 64'd0;
		mem_ctrl_memorycontroller836 <= 64'd0;
		mem_ctrl_memorycontroller837 <= 64'd0;
		mem_ctrl_memorycontroller838 <= 64'd0;
		mem_ctrl_memorycontroller839 <= 64'd0;
		mem_ctrl_memorycontroller840 <= 64'd0;
		mem_ctrl_memorycontroller841 <= 64'd0;
		mem_ctrl_memorycontroller842 <= 64'd0;
		mem_ctrl_memorycontroller843 <= 64'd0;
		mem_ctrl_memorycontroller844 <= 64'd0;
		mem_ctrl_memorycontroller845 <= 64'd0;
		mem_ctrl_memorycontroller846 <= 64'd0;
		mem_ctrl_memorycontroller847 <= 64'd0;
		mem_ctrl_memorycontroller848 <= 64'd0;
		mem_ctrl_memorycontroller849 <= 64'd0;
		mem_ctrl_memorycontroller850 <= 64'd0;
		mem_ctrl_memorycontroller851 <= 64'd0;
		mem_ctrl_memorycontroller852 <= 64'd0;
		mem_ctrl_memorycontroller853 <= 64'd0;
		mem_ctrl_memorycontroller854 <= 64'd0;
		mem_ctrl_memorycontroller855 <= 64'd0;
		mem_ctrl_memorycontroller856 <= 64'd0;
		mem_ctrl_memorycontroller857 <= 64'd0;
		mem_ctrl_memorycontroller858 <= 64'd0;
		mem_ctrl_memorycontroller859 <= 64'd0;
		mem_ctrl_memorycontroller860 <= 64'd0;
		mem_ctrl_memorycontroller861 <= 64'd0;
		mem_ctrl_memorycontroller862 <= 64'd0;
		mem_ctrl_memorycontroller863 <= 64'd0;
		mem_ctrl_memorycontroller864 <= 64'd0;
		mem_ctrl_memorycontroller865 <= 64'd0;
		mem_ctrl_memorycontroller866 <= 64'd0;
		mem_ctrl_memorycontroller867 <= 64'd0;
		mem_ctrl_memorycontroller868 <= 64'd0;
		mem_ctrl_memorycontroller869 <= 64'd0;
		mem_ctrl_memorycontroller870 <= 64'd0;
		mem_ctrl_memorycontroller871 <= 64'd0;
		mem_ctrl_memorycontroller872 <= 64'd0;
		mem_ctrl_memorycontroller873 <= 64'd0;
		mem_ctrl_memorycontroller874 <= 64'd0;
		mem_ctrl_memorycontroller875 <= 64'd0;
		mem_ctrl_memorycontroller876 <= 64'd0;
		mem_ctrl_memorycontroller877 <= 64'd0;
		mem_ctrl_memorycontroller878 <= 64'd0;
		mem_ctrl_memorycontroller879 <= 64'd0;
		mem_ctrl_memorycontroller880 <= 64'd0;
		mem_ctrl_memorycontroller881 <= 64'd0;
		mem_ctrl_memorycontroller882 <= 64'd0;
		mem_ctrl_memorycontroller883 <= 64'd0;
		mem_ctrl_memorycontroller884 <= 64'd0;
		mem_ctrl_memorycontroller885 <= 64'd0;
		mem_ctrl_memorycontroller886 <= 64'd0;
		mem_ctrl_memorycontroller887 <= 64'd0;
		mem_ctrl_memorycontroller888 <= 64'd0;
		mem_ctrl_memorycontroller889 <= 64'd0;
		mem_ctrl_memorycontroller890 <= 64'd0;
		mem_ctrl_memorycontroller891 <= 64'd0;
		mem_ctrl_memorycontroller892 <= 64'd0;
		mem_ctrl_memorycontroller893 <= 64'd0;
		mem_ctrl_memorycontroller894 <= 64'd0;
		mem_ctrl_memorycontroller895 <= 64'd0;
		mem_ctrl_memorycontroller896 <= 64'd0;
		mem_ctrl_memorycontroller897 <= 64'd0;
		mem_ctrl_memorycontroller898 <= 64'd0;
		mem_ctrl_memorycontroller899 <= 64'd0;
		mem_ctrl_memorycontroller900 <= 64'd0;
		mem_ctrl_memorycontroller901 <= 64'd0;
		mem_ctrl_memorycontroller902 <= 64'd0;
		mem_ctrl_memorycontroller903 <= 64'd0;
		mem_ctrl_memorycontroller904 <= 64'd0;
		mem_ctrl_memorycontroller905 <= 64'd0;
		mem_ctrl_memorycontroller906 <= 64'd0;
		mem_ctrl_memorycontroller907 <= 64'd0;
		mem_ctrl_memorycontroller908 <= 64'd0;
		mem_ctrl_memorycontroller909 <= 64'd0;
		mem_ctrl_memorycontroller910 <= 64'd0;
		mem_ctrl_memorycontroller911 <= 64'd0;
		mem_ctrl_memorycontroller912 <= 64'd0;
		mem_ctrl_memorycontroller913 <= 64'd0;
		mem_ctrl_memorycontroller914 <= 64'd0;
		mem_ctrl_memorycontroller915 <= 64'd0;
		mem_ctrl_memorycontroller916 <= 64'd0;
		mem_ctrl_memorycontroller917 <= 64'd0;
		mem_ctrl_memorycontroller918 <= 64'd0;
		mem_ctrl_memorycontroller919 <= 64'd0;
		mem_ctrl_memorycontroller920 <= 64'd0;
		mem_ctrl_memorycontroller921 <= 64'd0;
		mem_ctrl_memorycontroller922 <= 64'd0;
		mem_ctrl_memorycontroller923 <= 64'd0;
		mem_ctrl_memorycontroller924 <= 64'd0;
		mem_ctrl_memorycontroller925 <= 64'd0;
		mem_ctrl_memorycontroller926 <= 64'd0;
		mem_ctrl_memorycontroller927 <= 64'd0;
		mem_ctrl_memorycontroller928 <= 64'd0;
		mem_ctrl_memorycontroller929 <= 64'd0;
		mem_ctrl_memorycontroller930 <= 64'd0;
		mem_ctrl_memorycontroller931 <= 64'd0;
		mem_ctrl_memorycontroller932 <= 64'd0;
		mem_ctrl_memorycontroller933 <= 64'd0;
		mem_ctrl_memorycontroller934 <= 64'd0;
		mem_ctrl_memorycontroller935 <= 64'd0;
		mem_ctrl_memorycontroller936 <= 64'd0;
		mem_ctrl_memorycontroller937 <= 64'd0;
		mem_ctrl_memorycontroller938 <= 64'd0;
		mem_ctrl_memorycontroller939 <= 64'd0;
		mem_ctrl_memorycontroller940 <= 64'd0;
		mem_ctrl_memorycontroller941 <= 64'd0;
		mem_ctrl_memorycontroller942 <= 64'd0;
		mem_ctrl_memorycontroller943 <= 64'd0;
		mem_ctrl_memorycontroller944 <= 64'd0;
		mem_ctrl_memorycontroller945 <= 64'd0;
		mem_ctrl_memorycontroller946 <= 64'd0;
		mem_ctrl_memorycontroller947 <= 64'd0;
		mem_ctrl_memorycontroller948 <= 64'd0;
		mem_ctrl_memorycontroller949 <= 64'd0;
		mem_ctrl_memorycontroller950 <= 64'd0;
		mem_ctrl_memorycontroller951 <= 64'd0;
		mem_ctrl_memorycontroller952 <= 64'd0;
		mem_ctrl_memorycontroller953 <= 64'd0;
		mem_ctrl_memorycontroller954 <= 64'd0;
		mem_ctrl_memorycontroller955 <= 64'd0;
		mem_ctrl_memorycontroller956 <= 64'd0;
		mem_ctrl_memorycontroller957 <= 64'd0;
		mem_ctrl_memorycontroller958 <= 64'd0;
		mem_ctrl_memorycontroller959 <= 64'd0;
		mem_ctrl_memorycontroller960 <= 64'd0;
		mem_ctrl_memorycontroller961 <= 64'd0;
		mem_ctrl_memorycontroller962 <= 64'd0;
		mem_ctrl_memorycontroller963 <= 64'd0;
		mem_ctrl_memorycontroller964 <= 64'd0;
		mem_ctrl_memorycontroller965 <= 64'd0;
		mem_ctrl_memorycontroller966 <= 64'd0;
		mem_ctrl_memorycontroller967 <= 64'd0;
		mem_ctrl_memorycontroller968 <= 64'd0;
		mem_ctrl_memorycontroller969 <= 64'd0;
		mem_ctrl_memorycontroller970 <= 64'd0;
		mem_ctrl_memorycontroller971 <= 64'd0;
		mem_ctrl_memorycontroller972 <= 64'd0;
		mem_ctrl_memorycontroller973 <= 64'd0;
		mem_ctrl_memorycontroller974 <= 64'd0;
		mem_ctrl_memorycontroller975 <= 64'd0;
		mem_ctrl_memorycontroller976 <= 64'd0;
		mem_ctrl_memorycontroller977 <= 64'd0;
		mem_ctrl_memorycontroller978 <= 64'd0;
		mem_ctrl_memorycontroller979 <= 64'd0;
		mem_ctrl_memorycontroller980 <= 64'd0;
		mem_ctrl_memorycontroller981 <= 64'd0;
		mem_ctrl_memorycontroller982 <= 64'd0;
		mem_ctrl_memorycontroller983 <= 64'd0;
		mem_ctrl_memorycontroller984 <= 64'd0;
		mem_ctrl_memorycontroller985 <= 64'd0;
		mem_ctrl_memorycontroller986 <= 64'd0;
		mem_ctrl_memorycontroller987 <= 64'd0;
		mem_ctrl_memorycontroller988 <= 64'd0;
		mem_ctrl_memorycontroller989 <= 64'd0;
		mem_ctrl_memorycontroller990 <= 64'd0;
		mem_ctrl_memorycontroller991 <= 64'd0;
		mem_ctrl_memorycontroller992 <= 64'd0;
		mem_ctrl_memorycontroller993 <= 64'd0;
		mem_ctrl_memorycontroller994 <= 64'd0;
		mem_ctrl_memorycontroller995 <= 64'd0;
		mem_ctrl_memorycontroller996 <= 64'd0;
		mem_ctrl_memorycontroller997 <= 64'd0;
		mem_ctrl_memorycontroller998 <= 64'd0;
		mem_ctrl_memorycontroller999 <= 64'd0;
		mem_ctrl_memorycontroller1000 <= 64'd0;
		mem_ctrl_memorycontroller1001 <= 64'd0;
		mem_ctrl_memorycontroller1002 <= 64'd0;
		mem_ctrl_memorycontroller1003 <= 64'd0;
		mem_ctrl_memorycontroller1004 <= 64'd0;
		mem_ctrl_memorycontroller1005 <= 64'd0;
		mem_ctrl_memorycontroller1006 <= 64'd0;
		mem_ctrl_memorycontroller1007 <= 64'd0;
		mem_ctrl_memorycontroller1008 <= 64'd0;
		mem_ctrl_memorycontroller1009 <= 64'd0;
		mem_ctrl_memorycontroller1010 <= 64'd0;
		mem_ctrl_memorycontroller1011 <= 64'd0;
		mem_ctrl_memorycontroller1012 <= 64'd0;
		mem_ctrl_memorycontroller1013 <= 64'd0;
		mem_ctrl_memorycontroller1014 <= 64'd0;
		mem_ctrl_memorycontroller1015 <= 64'd0;
		mem_ctrl_memorycontroller1016 <= 64'd0;
		mem_ctrl_memorycontroller1017 <= 64'd0;
		mem_ctrl_memorycontroller1018 <= 64'd0;
		mem_ctrl_memorycontroller1019 <= 64'd0;
		mem_ctrl_memorycontroller1020 <= 64'd0;
		mem_ctrl_memorycontroller1021 <= 64'd0;
		mem_ctrl_memorycontroller1022 <= 64'd0;
		mem_ctrl_memorycontroller1023 <= 64'd0;
		mem_ctrl_memorycontroller1024 <= 64'd0;
		mem_ctrl_memorycontroller1025 <= 64'd0;
		mem_ctrl_memorycontroller1026 <= 64'd0;
		mem_ctrl_memorycontroller1027 <= 64'd0;
		mem_ctrl_memorycontroller1028 <= 64'd0;
		mem_ctrl_memorycontroller1029 <= 64'd0;
		mem_ctrl_memorycontroller1030 <= 64'd0;
		mem_ctrl_memorycontroller1031 <= 64'd0;
	end
end

endmodule
